module HardDrive(address,prog,dados_in,dados_out,write,clock,clock_a);
	input [31:0] address;
   input	[31:0] dados_in;
	input [31:0] prog;
	input clock, clock_a, write;
	output reg[31:0] dados_out;
	
	reg [31:0] HD[30719:0];
	
	initial begin
		//valores iniciais do hd
		
	
// programa zero: SO	
HD[0] = 32'b001101_11011_000000000000000000000; //['loadi', '$r27', '0']
HD[1] = 32'b001101_11101_000000000000000000000; //['loadi', '$r29', '0']
HD[2] = 32'b001101_11000_000000000000000000000; //['loadi', '$r24', '0']
HD[3] = 32'b001101_00000_000000000000000000000; //['loadi', '$r0', '0']
HD[4] = 32'b001101_11111_000000000000000000000; //['loadi', '$r31', '0']
HD[5] = 32'b001101_11010_000000000000000000000; //['loadi', '$r26', '0']
HD[6] = 32'b010000_00000_000000000000000000111; //['jmpi', 'main']
HD[7] = 32'b001101_00001_000000000000000000001; //['loadi', '$r1', '1']
HD[8] = 32'b001101_00011_000000000000000000001; //['loadi', '$r3', '1']
HD[9] = 32'b011011_00100_00001_00011_00000000000; //['eq', '$r4', '$r1', '$r3']
HD[10] = 32'b100010_00000_00100_0000011100000010; //['jei', '$r0', '$r4', 'L2']
HD[11] = 32'b001101_00011_000000000000000000100; //['loadi', '$r3', 4]
HD[12] = 32'b000001_00001_11000_00011_00000000000; //['add', '$r1', '$r24', '$r3']
HD[13] = 32'b001101_00100_000000000000000000000; //['loadi', '$r4', '0']
HD[14] = 32'b000001_00101_00001_00100_00000000000; //['add', '$r5', '$r1', '$r4']
HD[15] = 32'b001101_00001_000000000000000000000; //['loadi', '$r1', '0']
HD[16] = 32'b001110_00001_00101_0000000000000000; //['store', '$r1', '$r5']
HD[17] = 32'b001101_00011_000000000000000000100; //['loadi', '$r3', 4]
HD[18] = 32'b000001_00001_11000_00011_00000000000; //['add', '$r1', '$r24', '$r3']
HD[19] = 32'b001101_00100_000000000000000000001; //['loadi', '$r4', '1']
HD[20] = 32'b000001_00101_00001_00100_00000000000; //['add', '$r5', '$r1', '$r4']
HD[21] = 32'b001101_00001_000000000000000000000; //['loadi', '$r1', '0']
HD[22] = 32'b001110_00001_00101_0000000000000000; //['store', '$r1', '$r5']
HD[23] = 32'b001101_00011_000000000000000000100; //['loadi', '$r3', 4]
HD[24] = 32'b000001_00001_11000_00011_00000000000; //['add', '$r1', '$r24', '$r3']
HD[25] = 32'b001101_00100_000000000000000000010; //['loadi', '$r4', '2']
HD[26] = 32'b000001_00101_00001_00100_00000000000; //['add', '$r5', '$r1', '$r4']
HD[27] = 32'b001101_00001_000000000000000000000; //['loadi', '$r1', '0']
HD[28] = 32'b001110_00001_00101_0000000000000000; //['store', '$r1', '$r5']
HD[29] = 32'b001101_00011_000000000000000000100; //['loadi', '$r3', 4]
HD[30] = 32'b000001_00001_11000_00011_00000000000; //['add', '$r1', '$r24', '$r3']
HD[31] = 32'b001101_00100_000000000000000000011; //['loadi', '$r4', '3']
HD[32] = 32'b000001_00101_00001_00100_00000000000; //['add', '$r5', '$r1', '$r4']
HD[33] = 32'b001101_00001_000000000000000000000; //['loadi', '$r1', '0']
HD[34] = 32'b001110_00001_00101_0000000000000000; //['store', '$r1', '$r5']
HD[35] = 32'b001101_11110_000000000000000001111; //['loadi', '$r30', 15]
HD[36] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[37] = 32'b001101_00100_000000000000000000000; //['loadi', '$r4', '0']
HD[38] = 32'b001110_00100_00001_0000000000000000; //['store', '$r4', '$r1']
HD[39] = 32'b001101_11110_000000000000000010000; //['loadi', '$r30', 16]
HD[40] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[41] = 32'b001101_00100_000000000000000000000; //['loadi', '$r4', '0']
HD[42] = 32'b001110_00100_00001_0000000000000000; //['store', '$r4', '$r1']
HD[43] = 32'b001101_11110_000000000000000010001; //['loadi', '$r30', 17]
HD[44] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[45] = 32'b001101_00100_000000000000000000000; //['loadi', '$r4', '0']
HD[46] = 32'b001110_00100_00001_0000000000000000; //['store', '$r4', '$r1']
HD[47] = 32'b001101_11110_000000000000000010010; //['loadi', '$r30', 18]
HD[48] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[49] = 32'b001101_00100_000000000000000000000; //['loadi', '$r4', '0']
HD[50] = 32'b001110_00100_00001_0000000000000000; //['store', '$r4', '$r1']
HD[51] = 32'b001101_11110_000000000000000010011; //['loadi', '$r30', 19]
HD[52] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[53] = 32'b001101_00100_000000000000000000000; //['loadi', '$r4', '0']
HD[54] = 32'b001110_00100_00001_0000000000000000; //['store', '$r4', '$r1']
HD[55] = 32'b001101_11110_000000000000000010101; //['loadi', '$r30', 21]
HD[56] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[57] = 32'b001101_00100_000000000000000000001; //['loadi', '$r4', '1']
HD[58] = 32'b001110_00100_00001_0000000000000000; //['store', '$r4', '$r1']
HD[59] = 32'b001101_00011_000000000000000000000; //['loadi', '$r3', 0]
HD[60] = 32'b000001_00001_11000_00011_00000000000; //['add', '$r1', '$r24', '$r3']
HD[61] = 32'b001101_00100_000000000000000000000; //['loadi', '$r4', '0']
HD[62] = 32'b000001_00101_00001_00100_00000000000; //['add', '$r5', '$r1', '$r4']
HD[63] = 32'b001101_00001_000000000000000000000; //['loadi', '$r1', '0']
HD[64] = 32'b001110_00001_00101_0000000000000000; //['store', '$r1', '$r5']
HD[65] = 32'b001101_00011_000000000000000000000; //['loadi', '$r3', 0]
HD[66] = 32'b000001_00001_11000_00011_00000000000; //['add', '$r1', '$r24', '$r3']
HD[67] = 32'b001101_00100_000000000000000000001; //['loadi', '$r4', '1']
HD[68] = 32'b000001_00101_00001_00100_00000000000; //['add', '$r5', '$r1', '$r4']
HD[69] = 32'b001101_00001_000000000000000000000; //['loadi', '$r1', '0']
HD[70] = 32'b001110_00001_00101_0000000000000000; //['store', '$r1', '$r5']
HD[71] = 32'b001101_00011_000000000000000000000; //['loadi', '$r3', 0]
HD[72] = 32'b000001_00001_11000_00011_00000000000; //['add', '$r1', '$r24', '$r3']
HD[73] = 32'b001101_00100_000000000000000000010; //['loadi', '$r4', '2']
HD[74] = 32'b000001_00101_00001_00100_00000000000; //['add', '$r5', '$r1', '$r4']
HD[75] = 32'b001101_00001_000000000000000000000; //['loadi', '$r1', '0']
HD[76] = 32'b001110_00001_00101_0000000000000000; //['store', '$r1', '$r5']
HD[77] = 32'b001101_00011_000000000000000000000; //['loadi', '$r3', 0]
HD[78] = 32'b000001_00001_11000_00011_00000000000; //['add', '$r1', '$r24', '$r3']
HD[79] = 32'b001101_00100_000000000000000000011; //['loadi', '$r4', '3']
HD[80] = 32'b000001_00101_00001_00100_00000000000; //['add', '$r5', '$r1', '$r4']
HD[81] = 32'b001101_00001_000000000000000000000; //['loadi', '$r1', '0']
HD[82] = 32'b001110_00001_00101_0000000000000000; //['store', '$r1', '$r5']
HD[83] = 32'b001101_11110_000000000000000001110; //['loadi', '$r30', 14]
HD[84] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[85] = 32'b001101_00100_000000000000000000000; //['loadi', '$r4', '0']
HD[86] = 32'b001110_00100_00001_0000000000000000; //['store', '$r4', '$r1']
HD[87] = 32'b010110_11100_000000000000000000000; //['in', '$r28']
HD[88] = 32'b001111_00001_11100_0000000000000000; //['move', '$r1', '$r28']
HD[89] = 32'b001101_11110_000000000000000001101; //['loadi', '$r30', 13]
HD[90] = 32'b000001_00011_11000_11110_00000000000; //['add', '$r3', '$r24', '$r30']
HD[91] = 32'b001110_00001_00011_0000000000000000; //['store', '$r1', '$r3']
HD[92] = 32'b001101_11110_000000000000000001110; //['loadi', '$r30', 14]
HD[93] = 32'b000001_00011_11000_11110_00000000000; //['add', '$r3', '$r24', '$r30']
HD[94] = 32'b001100_00001_00011_0000000000000000; //['load', '$r1', '$r3']
HD[95] = 32'b001101_11110_000000000000000001101; //['loadi', '$r30', 13]
HD[96] = 32'b000001_00011_11000_11110_00000000000; //['add', '$r3', '$r24', '$r30']
HD[97] = 32'b001100_00100_00011_0000000000000000; //['load', '$r4', '$r3']
HD[98] = 32'b011111_00101_00001_00100_00000000000; //['lt', '$r5', '$r1', '$r4']
HD[99] = 32'b100010_00000_00101_0000000001110110; //['jei', '$r0', '$r5', 'L4']
HD[100] = 32'b010110_11100_000000000000000000000; //['in', '$r28']
HD[101] = 32'b001111_00001_11100_0000000000000000; //['move', '$r1', '$r28']
HD[102] = 32'b001101_00101_000000000000000000000; //['loadi', '$r5', 0]
HD[103] = 32'b000001_00100_11000_00101_00000000000; //['add', '$r4', '$r24', '$r5']
HD[104] = 32'b001101_11110_000000000000000001110; //['loadi', '$r30', 14]
HD[105] = 32'b000001_00101_11000_11110_00000000000; //['add', '$r5', '$r24', '$r30']
HD[106] = 32'b001100_00110_00101_0000000000000000; //['load', '$r6', '$r5']
HD[107] = 32'b000001_00111_00100_00110_00000000000; //['add', '$r7', '$r4', '$r6']
HD[108] = 32'b001110_00001_00111_0000000000000000; //['store', '$r1', '$r7']
HD[109] = 32'b001101_11110_000000000000000001110; //['loadi', '$r30', 14]
HD[110] = 32'b000001_00100_11000_11110_00000000000; //['add', '$r4', '$r24', '$r30']
HD[111] = 32'b001100_00001_00100_0000000000000000; //['load', '$r1', '$r4']
HD[112] = 32'b001101_00101_000000000000000000001; //['loadi', '$r5', '1']
HD[113] = 32'b000001_00110_00001_00101_00000000000; //['add', '$r6', '$r1', '$r5']
HD[114] = 32'b001101_11110_000000000000000001110; //['loadi', '$r30', 14]
HD[115] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[116] = 32'b001110_00110_00001_0000000000000000; //['store', '$r6', '$r1']
HD[117] = 32'b010000_00000_000000000000001011100; //['jmpi', 'L3']
HD[118] = 32'b001101_11110_000000000000000010011; //['loadi', '$r30', 19]
HD[119] = 32'b000001_00101_11000_11110_00000000000; //['add', '$r5', '$r24', '$r30']
HD[120] = 32'b001100_00001_00101_0000000000000000; //['load', '$r1', '$r5']
HD[121] = 32'b001101_11110_000000000000000001101; //['loadi', '$r30', 13]
HD[122] = 32'b000001_00101_11000_11110_00000000000; //['add', '$r5', '$r24', '$r30']
HD[123] = 32'b001100_00110_00101_0000000000000000; //['load', '$r6', '$r5']
HD[124] = 32'b011111_00111_00001_00110_00000000000; //['lt', '$r7', '$r1', '$r6']
HD[125] = 32'b100010_00000_00111_0000011100000001; //['jei', '$r0', '$r7', 'L6']
HD[126] = 32'b001101_00110_000000000000000000000; //['loadi', '$r6', 0]
HD[127] = 32'b000001_00001_11000_00110_00000000000; //['add', '$r1', '$r24', '$r6']
HD[128] = 32'b001101_11110_000000000000000010011; //['loadi', '$r30', 19]
HD[129] = 32'b000001_00110_11000_11110_00000000000; //['add', '$r6', '$r24', '$r30']
HD[130] = 32'b001100_00111_00110_0000000000000000; //['load', '$r7', '$r6']
HD[131] = 32'b000001_01001_00001_00111_00000000000; //['add', '$r9', '$r1', '$r7']
HD[132] = 32'b001100_01000_01001_0000000000000000; //['load', '$r8', '$r9']
HD[133] = 32'b001101_00001_000000000000000000000; //['loadi', '$r1', '0']
HD[134] = 32'b011101_00111_01000_00001_00000000000; //['abv', '$r7', '$r8', '$r1']
HD[135] = 32'b100010_00000_00111_0000011011000110; //['jei', '$r0', '$r7', 'L7']
HD[136] = 32'b001101_11110_000000000000000001000; //['loadi', '$r30', 8]
HD[137] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[138] = 32'b001101_01000_000000000000000000000; //['loadi', '$r8', '0']
HD[139] = 32'b001110_01000_00001_0000000000000000; //['store', '$r8', '$r1']
HD[140] = 32'b001101_11110_000000000000000001000; //['loadi', '$r30', 8]
HD[141] = 32'b000001_00111_11000_11110_00000000000; //['add', '$r7', '$r24', '$r30']
HD[142] = 32'b001100_00001_00111_0000000000000000; //['load', '$r1', '$r7']
HD[143] = 32'b001101_01000_000000000000001111000; //['loadi', '$r8', '120']
HD[144] = 32'b011111_01001_00001_01000_00000000000; //['lt', '$r9', '$r1', '$r8']
HD[145] = 32'b100010_00000_01001_0000000010101001; //['jei', '$r0', '$r9', 'L10']
HD[146] = 32'b001101_01000_000000000000000000000; //['loadi', '$r8', 0]
HD[147] = 32'b000001_00001_11000_01000_00000000000; //['add', '$r1', '$r24', '$r8']
HD[148] = 32'b001101_11110_000000000000000010011; //['loadi', '$r30', 19]
HD[149] = 32'b000001_01000_11000_11110_00000000000; //['add', '$r8', '$r24', '$r30']
HD[150] = 32'b001100_01001_01000_0000000000000000; //['load', '$r9', '$r8']
HD[151] = 32'b000001_01011_00001_01001_00000000000; //['add', '$r11', '$r1', '$r9']
HD[152] = 32'b001100_01010_01011_0000000000000000; //['load', '$r10', '$r11']
HD[153] = 32'b001101_11110_000000000000000001000; //['loadi', '$r30', 8]
HD[154] = 32'b000001_01000_11000_11110_00000000000; //['add', '$r8', '$r24', '$r30']
HD[155] = 32'b001100_00001_01000_0000000000000000; //['load', '$r1', '$r8']
HD[156] = 32'b001101_11110_000000000000000001000; //['loadi', '$r30', 8]
HD[157] = 32'b000001_01000_11000_11110_00000000000; //['add', '$r8', '$r24', '$r30']
HD[158] = 32'b001100_01001_01000_0000000000000000; //['load', '$r9', '$r8']
HD[159] = 32'b101001_01001_00001_01010_00000000000; //['movehdmem', '$r9', '$r1', '$r10']
HD[160] = 32'b001101_11110_000000000000000001000; //['loadi', '$r30', 8]
HD[161] = 32'b000001_01000_11000_11110_00000000000; //['add', '$r8', '$r24', '$r30']
HD[162] = 32'b001100_00001_01000_0000000000000000; //['load', '$r1', '$r8']
HD[163] = 32'b001101_01001_000000000000000000001; //['loadi', '$r9', '1']
HD[164] = 32'b000001_01010_00001_01001_00000000000; //['add', '$r10', '$r1', '$r9']
HD[165] = 32'b001101_11110_000000000000000001000; //['loadi', '$r30', 8]
HD[166] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[167] = 32'b001110_01010_00001_0000000000000000; //['store', '$r10', '$r1']
HD[168] = 32'b010000_00000_000000000000010001100; //['jmpi', 'L9']
HD[169] = 32'b001101_01001_000000000000000000100; //['loadi', '$r9', 4]
HD[170] = 32'b000001_00001_11000_01001_00000000000; //['add', '$r1', '$r24', '$r9']
HD[171] = 32'b001101_11110_000000000000000010011; //['loadi', '$r30', 19]
HD[172] = 32'b000001_01001_11000_11110_00000000000; //['add', '$r9', '$r24', '$r30']
HD[173] = 32'b001100_01010_01001_0000000000000000; //['load', '$r10', '$r9']
HD[174] = 32'b000001_01100_00001_01010_00000000000; //['add', '$r12', '$r1', '$r10']
HD[175] = 32'b001100_01011_01100_0000000000000000; //['load', '$r11', '$r12']
HD[176] = 32'b001101_00001_000000000000000000000; //['loadi', '$r1', '0']
HD[177] = 32'b011011_01010_01011_00001_00000000000; //['eq', '$r10', '$r11', '$r1']
HD[178] = 32'b100010_00000_01010_0000000011110000; //['jei', '$r0', '$r10', 'L11']
HD[179] = 32'b001101_11110_000000000000000010011; //['loadi', '$r30', 19]
HD[180] = 32'b000001_01010_11000_11110_00000000000; //['add', '$r10', '$r24', '$r30']
HD[181] = 32'b001100_00001_01010_0000000000000000; //['load', '$r1', '$r10']
HD[182] = 32'b001101_01011_000000000000000000000; //['loadi', '$r11', '0']
HD[183] = 32'b011011_01100_00001_01011_00000000000; //['eq', '$r12', '$r1', '$r11']
HD[184] = 32'b100010_00000_01100_0000000010111101; //['jei', '$r0', '$r12', 'L13']
HD[185] = 32'b001101_11110_000000000000000001001; //['loadi', '$r30', 9]
HD[186] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[187] = 32'b001101_01100_000000000001000000000; //['loadi', '$r12', '512']
HD[188] = 32'b001110_01100_00001_0000000000000000; //['store', '$r12', '$r1']
HD[189] = 32'b001101_11110_000000000000000010011; //['loadi', '$r30', 19]
HD[190] = 32'b000001_01011_11000_11110_00000000000; //['add', '$r11', '$r24', '$r30']
HD[191] = 32'b001100_00001_01011_0000000000000000; //['load', '$r1', '$r11']
HD[192] = 32'b001101_01100_000000000000000000001; //['loadi', '$r12', '1']
HD[193] = 32'b011011_01101_00001_01100_00000000000; //['eq', '$r13', '$r1', '$r12']
HD[194] = 32'b100010_00000_01101_0000000011000111; //['jei', '$r0', '$r13', 'L15']
HD[195] = 32'b001101_11110_000000000000000001001; //['loadi', '$r30', 9]
HD[196] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[197] = 32'b001101_01101_000000000010000000000; //['loadi', '$r13', '1024']
HD[198] = 32'b001110_01101_00001_0000000000000000; //['store', '$r13', '$r1']
HD[199] = 32'b001101_11110_000000000000000010011; //['loadi', '$r30', 19]
HD[200] = 32'b000001_01100_11000_11110_00000000000; //['add', '$r12', '$r24', '$r30']
HD[201] = 32'b001100_00001_01100_0000000000000000; //['load', '$r1', '$r12']
HD[202] = 32'b001101_01101_000000000000000000010; //['loadi', '$r13', '2']
HD[203] = 32'b011011_01110_00001_01101_00000000000; //['eq', '$r14', '$r1', '$r13']
HD[204] = 32'b100010_00000_01110_0000000011010001; //['jei', '$r0', '$r14', 'L17']
HD[205] = 32'b001101_11110_000000000000000001001; //['loadi', '$r30', 9]
HD[206] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[207] = 32'b001101_01110_000000000011000000000; //['loadi', '$r14', '1536']
HD[208] = 32'b001110_01110_00001_0000000000000000; //['store', '$r14', '$r1']
HD[209] = 32'b001101_11110_000000000000000010011; //['loadi', '$r30', 19]
HD[210] = 32'b000001_01101_11000_11110_00000000000; //['add', '$r13', '$r24', '$r30']
HD[211] = 32'b001100_00001_01101_0000000000000000; //['load', '$r1', '$r13']
HD[212] = 32'b001101_01110_000000000000000000011; //['loadi', '$r14', '3']
HD[213] = 32'b011011_01111_00001_01110_00000000000; //['eq', '$r15', '$r1', '$r14']
HD[214] = 32'b100010_00000_01111_0000000011011011; //['jei', '$r0', '$r15', 'L19']
HD[215] = 32'b001101_11110_000000000000000001001; //['loadi', '$r30', 9]
HD[216] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[217] = 32'b001101_01111_000000000100000000000; //['loadi', '$r15', '2048']
HD[218] = 32'b001110_01111_00001_0000000000000000; //['store', '$r15', '$r1']
HD[219] = 32'b001101_11110_000000000000000001001; //['loadi', '$r30', 9]
HD[220] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[221] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[222] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[223] = 32'b001111_11000_10110_0000000000000000; //['move', '$r24', '$r22']
HD[224] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[225] = 32'b001101_11110_000000000000000001001; //['loadi', '$r30', 9]
HD[226] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[227] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[228] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[229] = 32'b001111_11101_10110_0000000000000000; //['move', '$r29', '$r22']
HD[230] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[231] = 32'b001101_01110_000000000000000000100; //['loadi', '$r14', 4]
HD[232] = 32'b000001_00001_11000_01110_00000000000; //['add', '$r1', '$r24', '$r14']
HD[233] = 32'b001101_11110_000000000000000010011; //['loadi', '$r30', 19]
HD[234] = 32'b000001_01110_11000_11110_00000000000; //['add', '$r14', '$r24', '$r30']
HD[235] = 32'b001100_01111_01110_0000000000000000; //['load', '$r15', '$r14']
HD[236] = 32'b000001_10000_00001_01111_00000000000; //['add', '$r16', '$r1', '$r15']
HD[237] = 32'b001101_00001_000000000000000000001; //['loadi', '$r1', '1']
HD[238] = 32'b001110_00001_10000_0000000000000000; //['store', '$r1', '$r16']
HD[239] = 32'b010000_00000_000000000001110001000; //['jmpi', 'L12']
HD[240] = 32'b001101_11110_000000000000000010011; //['loadi', '$r30', 19]
HD[241] = 32'b000001_01110_11000_11110_00000000000; //['add', '$r14', '$r24', '$r30']
HD[242] = 32'b001100_00001_01110_0000000000000000; //['load', '$r1', '$r14']
HD[243] = 32'b001101_01111_000000000000000000000; //['loadi', '$r15', '0']
HD[244] = 32'b011011_10000_00001_01111_00000000000; //['eq', '$r16', '$r1', '$r15']
HD[245] = 32'b100010_00000_10000_0000000110010110; //['jei', '$r0', '$r16', 'L21']
HD[246] = 32'b001101_00001_000000000000110010000; //['loadi', '$r1', '400']
HD[247] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[248] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[249] = 32'b001111_00000_10110_0000000000000000; //['move', '$r0', '$r22']
HD[250] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[251] = 32'b001101_00001_000000000000110010001; //['loadi', '$r1', '401']
HD[252] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[253] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[254] = 32'b001111_00001_10110_0000000000000000; //['move', '$r1', '$r22']
HD[255] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[256] = 32'b001101_00001_000000000000110010010; //['loadi', '$r1', '402']
HD[257] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[258] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[259] = 32'b001111_00010_10110_0000000000000000; //['move', '$r2', '$r22']
HD[260] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[261] = 32'b001101_00001_000000000000110010011; //['loadi', '$r1', '403']
HD[262] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[263] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[264] = 32'b001111_00011_10110_0000000000000000; //['move', '$r3', '$r22']
HD[265] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[266] = 32'b001101_00001_000000000000110010100; //['loadi', '$r1', '404']
HD[267] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[268] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[269] = 32'b001111_00100_10110_0000000000000000; //['move', '$r4', '$r22']
HD[270] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[271] = 32'b001101_00001_000000000000110010101; //['loadi', '$r1', '405']
HD[272] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[273] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[274] = 32'b001111_00101_10110_0000000000000000; //['move', '$r5', '$r22']
HD[275] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[276] = 32'b001101_00001_000000000000110010110; //['loadi', '$r1', '406']
HD[277] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[278] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[279] = 32'b001111_00110_10110_0000000000000000; //['move', '$r6', '$r22']
HD[280] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[281] = 32'b001101_00001_000000000000110010111; //['loadi', '$r1', '407']
HD[282] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[283] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[284] = 32'b001111_00111_10110_0000000000000000; //['move', '$r7', '$r22']
HD[285] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[286] = 32'b001101_00001_000000000000110011000; //['loadi', '$r1', '408']
HD[287] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[288] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[289] = 32'b001111_01000_10110_0000000000000000; //['move', '$r8', '$r22']
HD[290] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[291] = 32'b001101_00001_000000000000110011001; //['loadi', '$r1', '409']
HD[292] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[293] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[294] = 32'b001111_01001_10110_0000000000000000; //['move', '$r9', '$r22']
HD[295] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[296] = 32'b001101_00001_000000000000110011010; //['loadi', '$r1', '410']
HD[297] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[298] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[299] = 32'b001111_01010_10110_0000000000000000; //['move', '$r10', '$r22']
HD[300] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[301] = 32'b001101_00001_000000000000110011011; //['loadi', '$r1', '411']
HD[302] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[303] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[304] = 32'b001111_01011_10110_0000000000000000; //['move', '$r11', '$r22']
HD[305] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[306] = 32'b001101_00001_000000000000110011100; //['loadi', '$r1', '412']
HD[307] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[308] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[309] = 32'b001111_01100_10110_0000000000000000; //['move', '$r12', '$r22']
HD[310] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[311] = 32'b001101_00001_000000000000110011101; //['loadi', '$r1', '413']
HD[312] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[313] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[314] = 32'b001111_01101_10110_0000000000000000; //['move', '$r13', '$r22']
HD[315] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[316] = 32'b001101_00001_000000000000110011110; //['loadi', '$r1', '414']
HD[317] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[318] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[319] = 32'b001111_01110_10110_0000000000000000; //['move', '$r14', '$r22']
HD[320] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[321] = 32'b001101_00001_000000000000110011111; //['loadi', '$r1', '415']
HD[322] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[323] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[324] = 32'b001111_01111_10110_0000000000000000; //['move', '$r15', '$r22']
HD[325] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[326] = 32'b001101_00001_000000000000110100000; //['loadi', '$r1', '416']
HD[327] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[328] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[329] = 32'b001111_10000_10110_0000000000000000; //['move', '$r16', '$r22']
HD[330] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[331] = 32'b001101_00001_000000000000110100001; //['loadi', '$r1', '417']
HD[332] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[333] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[334] = 32'b001111_10001_10110_0000000000000000; //['move', '$r17', '$r22']
HD[335] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[336] = 32'b001101_00001_000000000000110100010; //['loadi', '$r1', '418']
HD[337] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[338] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[339] = 32'b001111_10010_10110_0000000000000000; //['move', '$r18', '$r22']
HD[340] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[341] = 32'b001101_00001_000000000000110100011; //['loadi', '$r1', '419']
HD[342] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[343] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[344] = 32'b001111_10011_10110_0000000000000000; //['move', '$r19', '$r22']
HD[345] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[346] = 32'b001101_00001_000000000000110100100; //['loadi', '$r1', '420']
HD[347] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[348] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[349] = 32'b001111_10100_10110_0000000000000000; //['move', '$r20', '$r22']
HD[350] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[351] = 32'b001101_00001_000000000000110100101; //['loadi', '$r1', '421']
HD[352] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[353] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[354] = 32'b001111_10101_10110_0000000000000000; //['move', '$r21', '$r22']
HD[355] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[356] = 32'b001101_00001_000000000000110100110; //['loadi', '$r1', '422']
HD[357] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[358] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[359] = 32'b001111_10110_10110_0000000000000000; //['move', '$r22', '$r22']
HD[360] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[361] = 32'b001101_00001_000000000000110100111; //['loadi', '$r1', '423']
HD[362] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[363] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[364] = 32'b001111_10111_10110_0000000000000000; //['move', '$r23', '$r22']
HD[365] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[366] = 32'b001101_00001_000000000000110101000; //['loadi', '$r1', '424']
HD[367] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[368] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[369] = 32'b001111_11000_10110_0000000000000000; //['move', '$r24', '$r22']
HD[370] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[371] = 32'b001101_00001_000000000000110101001; //['loadi', '$r1', '425']
HD[372] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[373] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[374] = 32'b001111_11001_10110_0000000000000000; //['move', '$r25', '$r22']
HD[375] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[376] = 32'b001101_00001_000000000000110101010; //['loadi', '$r1', '426']
HD[377] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[378] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[379] = 32'b001111_11010_10110_0000000000000000; //['move', '$r26', '$r22']
HD[380] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[381] = 32'b001101_00001_000000000000110101011; //['loadi', '$r1', '427']
HD[382] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[383] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[384] = 32'b001111_11011_10110_0000000000000000; //['move', '$r27', '$r22']
HD[385] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[386] = 32'b001101_00001_000000000000110101100; //['loadi', '$r1', '428']
HD[387] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[388] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[389] = 32'b001111_11100_10110_0000000000000000; //['move', '$r28', '$r22']
HD[390] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[391] = 32'b001101_00001_000000000000110101101; //['loadi', '$r1', '429']
HD[392] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[393] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[394] = 32'b001111_11101_10110_0000000000000000; //['move', '$r29', '$r22']
HD[395] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[396] = 32'b001101_00001_000000000000110101110; //['loadi', '$r1', '430']
HD[397] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[398] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[399] = 32'b001111_11110_10110_0000000000000000; //['move', '$r30', '$r22']
HD[400] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[401] = 32'b001101_00001_000000000000110101111; //['loadi', '$r1', '431']
HD[402] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[403] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[404] = 32'b001111_11111_10110_0000000000000000; //['move', '$r31', '$r22']
HD[405] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[406] = 32'b001101_11110_000000000000000010011; //['loadi', '$r30', 19]
HD[407] = 32'b000001_01111_11000_11110_00000000000; //['add', '$r15', '$r24', '$r30']
HD[408] = 32'b001100_00001_01111_0000000000000000; //['load', '$r1', '$r15']
HD[409] = 32'b001101_10000_000000000000000000001; //['loadi', '$r16', '1']
HD[410] = 32'b011011_10001_00001_10000_00000000000; //['eq', '$r17', '$r1', '$r16']
HD[411] = 32'b100010_00000_10001_0000001000111100; //['jei', '$r0', '$r17', 'L23']
HD[412] = 32'b001101_00001_000000000000110110000; //['loadi', '$r1', '432']
HD[413] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[414] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[415] = 32'b001111_00000_10110_0000000000000000; //['move', '$r0', '$r22']
HD[416] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[417] = 32'b001101_00001_000000000000110110001; //['loadi', '$r1', '433']
HD[418] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[419] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[420] = 32'b001111_00001_10110_0000000000000000; //['move', '$r1', '$r22']
HD[421] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[422] = 32'b001101_00001_000000000000110110010; //['loadi', '$r1', '434']
HD[423] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[424] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[425] = 32'b001111_00010_10110_0000000000000000; //['move', '$r2', '$r22']
HD[426] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[427] = 32'b001101_00001_000000000000110110011; //['loadi', '$r1', '435']
HD[428] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[429] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[430] = 32'b001111_00011_10110_0000000000000000; //['move', '$r3', '$r22']
HD[431] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[432] = 32'b001101_00001_000000000000110110100; //['loadi', '$r1', '436']
HD[433] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[434] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[435] = 32'b001111_00100_10110_0000000000000000; //['move', '$r4', '$r22']
HD[436] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[437] = 32'b001101_00001_000000000000110110101; //['loadi', '$r1', '437']
HD[438] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[439] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[440] = 32'b001111_00101_10110_0000000000000000; //['move', '$r5', '$r22']
HD[441] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[442] = 32'b001101_00001_000000000000110110110; //['loadi', '$r1', '438']
HD[443] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[444] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[445] = 32'b001111_00110_10110_0000000000000000; //['move', '$r6', '$r22']
HD[446] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[447] = 32'b001101_00001_000000000000110110111; //['loadi', '$r1', '439']
HD[448] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[449] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[450] = 32'b001111_00111_10110_0000000000000000; //['move', '$r7', '$r22']
HD[451] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[452] = 32'b001101_00001_000000000000110111000; //['loadi', '$r1', '440']
HD[453] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[454] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[455] = 32'b001111_01000_10110_0000000000000000; //['move', '$r8', '$r22']
HD[456] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[457] = 32'b001101_00001_000000000000110111001; //['loadi', '$r1', '441']
HD[458] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[459] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[460] = 32'b001111_01001_10110_0000000000000000; //['move', '$r9', '$r22']
HD[461] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[462] = 32'b001101_00001_000000000000110111010; //['loadi', '$r1', '442']
HD[463] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[464] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[465] = 32'b001111_01010_10110_0000000000000000; //['move', '$r10', '$r22']
HD[466] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[467] = 32'b001101_00001_000000000000110111011; //['loadi', '$r1', '443']
HD[468] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[469] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[470] = 32'b001111_01011_10110_0000000000000000; //['move', '$r11', '$r22']
HD[471] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[472] = 32'b001101_00001_000000000000110111100; //['loadi', '$r1', '444']
HD[473] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[474] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[475] = 32'b001111_01100_10110_0000000000000000; //['move', '$r12', '$r22']
HD[476] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[477] = 32'b001101_00001_000000000000110111101; //['loadi', '$r1', '445']
HD[478] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[479] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[480] = 32'b001111_01101_10110_0000000000000000; //['move', '$r13', '$r22']
HD[481] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[482] = 32'b001101_00001_000000000000110111110; //['loadi', '$r1', '446']
HD[483] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[484] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[485] = 32'b001111_01110_10110_0000000000000000; //['move', '$r14', '$r22']
HD[486] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[487] = 32'b001101_00001_000000000000110111111; //['loadi', '$r1', '447']
HD[488] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[489] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[490] = 32'b001111_01111_10110_0000000000000000; //['move', '$r15', '$r22']
HD[491] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[492] = 32'b001101_00001_000000000000111000000; //['loadi', '$r1', '448']
HD[493] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[494] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[495] = 32'b001111_10000_10110_0000000000000000; //['move', '$r16', '$r22']
HD[496] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[497] = 32'b001101_00001_000000000000111000001; //['loadi', '$r1', '449']
HD[498] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[499] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[500] = 32'b001111_10001_10110_0000000000000000; //['move', '$r17', '$r22']
HD[501] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[502] = 32'b001101_00001_000000000000111000010; //['loadi', '$r1', '450']
HD[503] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[504] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[505] = 32'b001111_10010_10110_0000000000000000; //['move', '$r18', '$r22']
HD[506] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[507] = 32'b001101_00001_000000000000111000011; //['loadi', '$r1', '451']
HD[508] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[509] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[510] = 32'b001111_10011_10110_0000000000000000; //['move', '$r19', '$r22']
HD[511] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[512] = 32'b001101_00001_000000000000111000100; //['loadi', '$r1', '452']
HD[513] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[514] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[515] = 32'b001111_10100_10110_0000000000000000; //['move', '$r20', '$r22']
HD[516] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[517] = 32'b001101_00001_000000000000111000101; //['loadi', '$r1', '453']
HD[518] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[519] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[520] = 32'b001111_10101_10110_0000000000000000; //['move', '$r21', '$r22']
HD[521] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[522] = 32'b001101_00001_000000000000111000110; //['loadi', '$r1', '454']
HD[523] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[524] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[525] = 32'b001111_10110_10110_0000000000000000; //['move', '$r22', '$r22']
HD[526] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[527] = 32'b001101_00001_000000000000111000111; //['loadi', '$r1', '455']
HD[528] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[529] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[530] = 32'b001111_10111_10110_0000000000000000; //['move', '$r23', '$r22']
HD[531] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[532] = 32'b001101_00001_000000000000111001000; //['loadi', '$r1', '456']
HD[533] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[534] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[535] = 32'b001111_11000_10110_0000000000000000; //['move', '$r24', '$r22']
HD[536] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[537] = 32'b001101_00001_000000000000111001001; //['loadi', '$r1', '457']
HD[538] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[539] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[540] = 32'b001111_11001_10110_0000000000000000; //['move', '$r25', '$r22']
HD[541] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[542] = 32'b001101_00001_000000000000111001010; //['loadi', '$r1', '458']
HD[543] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[544] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[545] = 32'b001111_11010_10110_0000000000000000; //['move', '$r26', '$r22']
HD[546] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[547] = 32'b001101_00001_000000000000111001011; //['loadi', '$r1', '459']
HD[548] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[549] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[550] = 32'b001111_11011_10110_0000000000000000; //['move', '$r27', '$r22']
HD[551] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[552] = 32'b001101_00001_000000000000111001100; //['loadi', '$r1', '460']
HD[553] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[554] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[555] = 32'b001111_11100_10110_0000000000000000; //['move', '$r28', '$r22']
HD[556] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[557] = 32'b001101_00001_000000000000111001101; //['loadi', '$r1', '461']
HD[558] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[559] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[560] = 32'b001111_11101_10110_0000000000000000; //['move', '$r29', '$r22']
HD[561] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[562] = 32'b001101_00001_000000000000111001110; //['loadi', '$r1', '462']
HD[563] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[564] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[565] = 32'b001111_11110_10110_0000000000000000; //['move', '$r30', '$r22']
HD[566] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[567] = 32'b001101_00001_000000000000111001111; //['loadi', '$r1', '463']
HD[568] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[569] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[570] = 32'b001111_11111_10110_0000000000000000; //['move', '$r31', '$r22']
HD[571] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[572] = 32'b001101_11110_000000000000000010011; //['loadi', '$r30', 19]
HD[573] = 32'b000001_10000_11000_11110_00000000000; //['add', '$r16', '$r24', '$r30']
HD[574] = 32'b001100_00001_10000_0000000000000000; //['load', '$r1', '$r16']
HD[575] = 32'b001101_10001_000000000000000000010; //['loadi', '$r17', '2']
HD[576] = 32'b011011_10010_00001_10001_00000000000; //['eq', '$r18', '$r1', '$r17']
HD[577] = 32'b100010_00000_10010_0000001011100010; //['jei', '$r0', '$r18', 'L25']
HD[578] = 32'b001101_00001_000000000000100101100; //['loadi', '$r1', '300']
HD[579] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[580] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[581] = 32'b001111_00000_10110_0000000000000000; //['move', '$r0', '$r22']
HD[582] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[583] = 32'b001101_00001_000000000000100101101; //['loadi', '$r1', '301']
HD[584] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[585] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[586] = 32'b001111_00001_10110_0000000000000000; //['move', '$r1', '$r22']
HD[587] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[588] = 32'b001101_00001_000000000000100101110; //['loadi', '$r1', '302']
HD[589] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[590] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[591] = 32'b001111_00010_10110_0000000000000000; //['move', '$r2', '$r22']
HD[592] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[593] = 32'b001101_00001_000000000000100101111; //['loadi', '$r1', '303']
HD[594] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[595] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[596] = 32'b001111_00011_10110_0000000000000000; //['move', '$r3', '$r22']
HD[597] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[598] = 32'b001101_00001_000000000000100110000; //['loadi', '$r1', '304']
HD[599] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[600] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[601] = 32'b001111_00100_10110_0000000000000000; //['move', '$r4', '$r22']
HD[602] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[603] = 32'b001101_00001_000000000000100110001; //['loadi', '$r1', '305']
HD[604] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[605] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[606] = 32'b001111_00101_10110_0000000000000000; //['move', '$r5', '$r22']
HD[607] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[608] = 32'b001101_00001_000000000000100110010; //['loadi', '$r1', '306']
HD[609] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[610] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[611] = 32'b001111_00110_10110_0000000000000000; //['move', '$r6', '$r22']
HD[612] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[613] = 32'b001101_00001_000000000000100110011; //['loadi', '$r1', '307']
HD[614] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[615] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[616] = 32'b001111_00111_10110_0000000000000000; //['move', '$r7', '$r22']
HD[617] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[618] = 32'b001101_00001_000000000000100110100; //['loadi', '$r1', '308']
HD[619] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[620] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[621] = 32'b001111_01000_10110_0000000000000000; //['move', '$r8', '$r22']
HD[622] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[623] = 32'b001101_00001_000000000000100110101; //['loadi', '$r1', '309']
HD[624] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[625] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[626] = 32'b001111_01001_10110_0000000000000000; //['move', '$r9', '$r22']
HD[627] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[628] = 32'b001101_00001_000000000000100110110; //['loadi', '$r1', '310']
HD[629] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[630] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[631] = 32'b001111_01010_10110_0000000000000000; //['move', '$r10', '$r22']
HD[632] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[633] = 32'b001101_00001_000000000000100110111; //['loadi', '$r1', '311']
HD[634] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[635] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[636] = 32'b001111_01011_10110_0000000000000000; //['move', '$r11', '$r22']
HD[637] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[638] = 32'b001101_00001_000000000000100111000; //['loadi', '$r1', '312']
HD[639] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[640] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[641] = 32'b001111_01100_10110_0000000000000000; //['move', '$r12', '$r22']
HD[642] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[643] = 32'b001101_00001_000000000000100111001; //['loadi', '$r1', '313']
HD[644] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[645] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[646] = 32'b001111_01101_10110_0000000000000000; //['move', '$r13', '$r22']
HD[647] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[648] = 32'b001101_00001_000000000000100111010; //['loadi', '$r1', '314']
HD[649] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[650] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[651] = 32'b001111_01110_10110_0000000000000000; //['move', '$r14', '$r22']
HD[652] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[653] = 32'b001101_00001_000000000000100111011; //['loadi', '$r1', '315']
HD[654] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[655] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[656] = 32'b001111_01111_10110_0000000000000000; //['move', '$r15', '$r22']
HD[657] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[658] = 32'b001101_00001_000000000000100111100; //['loadi', '$r1', '316']
HD[659] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[660] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[661] = 32'b001111_10000_10110_0000000000000000; //['move', '$r16', '$r22']
HD[662] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[663] = 32'b001101_00001_000000000000100111101; //['loadi', '$r1', '317']
HD[664] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[665] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[666] = 32'b001111_10001_10110_0000000000000000; //['move', '$r17', '$r22']
HD[667] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[668] = 32'b001101_00001_000000000000100111110; //['loadi', '$r1', '318']
HD[669] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[670] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[671] = 32'b001111_10010_10110_0000000000000000; //['move', '$r18', '$r22']
HD[672] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[673] = 32'b001101_00001_000000000000100111111; //['loadi', '$r1', '319']
HD[674] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[675] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[676] = 32'b001111_10011_10110_0000000000000000; //['move', '$r19', '$r22']
HD[677] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[678] = 32'b001101_00001_000000000000101000000; //['loadi', '$r1', '320']
HD[679] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[680] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[681] = 32'b001111_10100_10110_0000000000000000; //['move', '$r20', '$r22']
HD[682] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[683] = 32'b001101_00001_000000000000101000001; //['loadi', '$r1', '321']
HD[684] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[685] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[686] = 32'b001111_10101_10110_0000000000000000; //['move', '$r21', '$r22']
HD[687] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[688] = 32'b001101_00001_000000000000101000010; //['loadi', '$r1', '322']
HD[689] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[690] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[691] = 32'b001111_10110_10110_0000000000000000; //['move', '$r22', '$r22']
HD[692] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[693] = 32'b001101_00001_000000000000101000011; //['loadi', '$r1', '323']
HD[694] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[695] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[696] = 32'b001111_10111_10110_0000000000000000; //['move', '$r23', '$r22']
HD[697] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[698] = 32'b001101_00001_000000000000101000100; //['loadi', '$r1', '324']
HD[699] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[700] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[701] = 32'b001111_11000_10110_0000000000000000; //['move', '$r24', '$r22']
HD[702] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[703] = 32'b001101_00001_000000000000101000101; //['loadi', '$r1', '325']
HD[704] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[705] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[706] = 32'b001111_11001_10110_0000000000000000; //['move', '$r25', '$r22']
HD[707] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[708] = 32'b001101_00001_000000000000101000110; //['loadi', '$r1', '326']
HD[709] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[710] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[711] = 32'b001111_11010_10110_0000000000000000; //['move', '$r26', '$r22']
HD[712] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[713] = 32'b001101_00001_000000000000101000111; //['loadi', '$r1', '327']
HD[714] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[715] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[716] = 32'b001111_11011_10110_0000000000000000; //['move', '$r27', '$r22']
HD[717] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[718] = 32'b001101_00001_000000000000101001000; //['loadi', '$r1', '328']
HD[719] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[720] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[721] = 32'b001111_11100_10110_0000000000000000; //['move', '$r28', '$r22']
HD[722] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[723] = 32'b001101_00001_000000000000101001001; //['loadi', '$r1', '329']
HD[724] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[725] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[726] = 32'b001111_11101_10110_0000000000000000; //['move', '$r29', '$r22']
HD[727] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[728] = 32'b001101_00001_000000000000101001010; //['loadi', '$r1', '330']
HD[729] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[730] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[731] = 32'b001111_11110_10110_0000000000000000; //['move', '$r30', '$r22']
HD[732] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[733] = 32'b001101_00001_000000000000101001011; //['loadi', '$r1', '331']
HD[734] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[735] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[736] = 32'b001111_11111_10110_0000000000000000; //['move', '$r31', '$r22']
HD[737] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[738] = 32'b001101_11110_000000000000000010011; //['loadi', '$r30', 19]
HD[739] = 32'b000001_10001_11000_11110_00000000000; //['add', '$r17', '$r24', '$r30']
HD[740] = 32'b001100_00001_10001_0000000000000000; //['load', '$r1', '$r17']
HD[741] = 32'b001101_10010_000000000000000000011; //['loadi', '$r18', '3']
HD[742] = 32'b011011_10011_00001_10010_00000000000; //['eq', '$r19', '$r1', '$r18']
HD[743] = 32'b100010_00000_10011_0000001110001000; //['jei', '$r0', '$r19', 'L27']
HD[744] = 32'b001101_00001_000000000000101001100; //['loadi', '$r1', '332']
HD[745] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[746] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[747] = 32'b001111_00000_10110_0000000000000000; //['move', '$r0', '$r22']
HD[748] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[749] = 32'b001101_00001_000000000000101001101; //['loadi', '$r1', '333']
HD[750] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[751] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[752] = 32'b001111_00001_10110_0000000000000000; //['move', '$r1', '$r22']
HD[753] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[754] = 32'b001101_00001_000000000000101001110; //['loadi', '$r1', '334']
HD[755] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[756] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[757] = 32'b001111_00010_10110_0000000000000000; //['move', '$r2', '$r22']
HD[758] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[759] = 32'b001101_00001_000000000000101001111; //['loadi', '$r1', '335']
HD[760] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[761] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[762] = 32'b001111_00011_10110_0000000000000000; //['move', '$r3', '$r22']
HD[763] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[764] = 32'b001101_00001_000000000000101010000; //['loadi', '$r1', '336']
HD[765] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[766] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[767] = 32'b001111_00100_10110_0000000000000000; //['move', '$r4', '$r22']
HD[768] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[769] = 32'b001101_00001_000000000000101010001; //['loadi', '$r1', '337']
HD[770] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[771] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[772] = 32'b001111_00101_10110_0000000000000000; //['move', '$r5', '$r22']
HD[773] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[774] = 32'b001101_00001_000000000000101010010; //['loadi', '$r1', '338']
HD[775] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[776] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[777] = 32'b001111_00110_10110_0000000000000000; //['move', '$r6', '$r22']
HD[778] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[779] = 32'b001101_00001_000000000000101010011; //['loadi', '$r1', '339']
HD[780] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[781] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[782] = 32'b001111_00111_10110_0000000000000000; //['move', '$r7', '$r22']
HD[783] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[784] = 32'b001101_00001_000000000000101010100; //['loadi', '$r1', '340']
HD[785] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[786] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[787] = 32'b001111_01000_10110_0000000000000000; //['move', '$r8', '$r22']
HD[788] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[789] = 32'b001101_00001_000000000000101010101; //['loadi', '$r1', '341']
HD[790] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[791] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[792] = 32'b001111_01001_10110_0000000000000000; //['move', '$r9', '$r22']
HD[793] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[794] = 32'b001101_00001_000000000000101010110; //['loadi', '$r1', '342']
HD[795] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[796] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[797] = 32'b001111_01010_10110_0000000000000000; //['move', '$r10', '$r22']
HD[798] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[799] = 32'b001101_00001_000000000000101010111; //['loadi', '$r1', '343']
HD[800] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[801] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[802] = 32'b001111_01011_10110_0000000000000000; //['move', '$r11', '$r22']
HD[803] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[804] = 32'b001101_00001_000000000000101011000; //['loadi', '$r1', '344']
HD[805] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[806] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[807] = 32'b001111_01100_10110_0000000000000000; //['move', '$r12', '$r22']
HD[808] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[809] = 32'b001101_00001_000000000000101011001; //['loadi', '$r1', '345']
HD[810] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[811] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[812] = 32'b001111_01101_10110_0000000000000000; //['move', '$r13', '$r22']
HD[813] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[814] = 32'b001101_00001_000000000000101011010; //['loadi', '$r1', '346']
HD[815] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[816] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[817] = 32'b001111_01110_10110_0000000000000000; //['move', '$r14', '$r22']
HD[818] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[819] = 32'b001101_00001_000000000000101011011; //['loadi', '$r1', '347']
HD[820] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[821] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[822] = 32'b001111_01111_10110_0000000000000000; //['move', '$r15', '$r22']
HD[823] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[824] = 32'b001101_00001_000000000000101011100; //['loadi', '$r1', '348']
HD[825] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[826] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[827] = 32'b001111_10000_10110_0000000000000000; //['move', '$r16', '$r22']
HD[828] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[829] = 32'b001101_00001_000000000000101011101; //['loadi', '$r1', '349']
HD[830] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[831] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[832] = 32'b001111_10001_10110_0000000000000000; //['move', '$r17', '$r22']
HD[833] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[834] = 32'b001101_00001_000000000000101011110; //['loadi', '$r1', '350']
HD[835] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[836] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[837] = 32'b001111_10010_10110_0000000000000000; //['move', '$r18', '$r22']
HD[838] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[839] = 32'b001101_00001_000000000000101011111; //['loadi', '$r1', '351']
HD[840] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[841] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[842] = 32'b001111_10011_10110_0000000000000000; //['move', '$r19', '$r22']
HD[843] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[844] = 32'b001101_00001_000000000000101100000; //['loadi', '$r1', '352']
HD[845] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[846] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[847] = 32'b001111_10100_10110_0000000000000000; //['move', '$r20', '$r22']
HD[848] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[849] = 32'b001101_00001_000000000000101100001; //['loadi', '$r1', '353']
HD[850] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[851] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[852] = 32'b001111_10101_10110_0000000000000000; //['move', '$r21', '$r22']
HD[853] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[854] = 32'b001101_00001_000000000000101100010; //['loadi', '$r1', '354']
HD[855] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[856] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[857] = 32'b001111_10110_10110_0000000000000000; //['move', '$r22', '$r22']
HD[858] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[859] = 32'b001101_00001_000000000000101100011; //['loadi', '$r1', '355']
HD[860] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[861] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[862] = 32'b001111_10111_10110_0000000000000000; //['move', '$r23', '$r22']
HD[863] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[864] = 32'b001101_00001_000000000000101100100; //['loadi', '$r1', '356']
HD[865] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[866] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[867] = 32'b001111_11000_10110_0000000000000000; //['move', '$r24', '$r22']
HD[868] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[869] = 32'b001101_00001_000000000000101100101; //['loadi', '$r1', '357']
HD[870] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[871] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[872] = 32'b001111_11001_10110_0000000000000000; //['move', '$r25', '$r22']
HD[873] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[874] = 32'b001101_00001_000000000000101100110; //['loadi', '$r1', '358']
HD[875] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[876] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[877] = 32'b001111_11010_10110_0000000000000000; //['move', '$r26', '$r22']
HD[878] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[879] = 32'b001101_00001_000000000000101100111; //['loadi', '$r1', '359']
HD[880] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[881] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[882] = 32'b001111_11011_10110_0000000000000000; //['move', '$r27', '$r22']
HD[883] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[884] = 32'b001101_00001_000000000000101101000; //['loadi', '$r1', '360']
HD[885] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[886] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[887] = 32'b001111_11100_10110_0000000000000000; //['move', '$r28', '$r22']
HD[888] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[889] = 32'b001101_00001_000000000000101101001; //['loadi', '$r1', '361']
HD[890] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[891] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[892] = 32'b001111_11101_10110_0000000000000000; //['move', '$r29', '$r22']
HD[893] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[894] = 32'b001101_00001_000000000000101101010; //['loadi', '$r1', '362']
HD[895] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[896] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[897] = 32'b001111_11110_10110_0000000000000000; //['move', '$r30', '$r22']
HD[898] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[899] = 32'b001101_00001_000000000000101101011; //['loadi', '$r1', '363']
HD[900] = 32'b001100_10110_00001_0000000000000000; //['load', '$r22', '$r1']
HD[901] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[902] = 32'b001111_11111_10110_0000000000000000; //['move', '$r31', '$r22']
HD[903] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[904] = 32'b001101_11110_000000000000000010011; //['loadi', '$r30', 19]
HD[905] = 32'b000001_10010_11000_11110_00000000000; //['add', '$r18', '$r24', '$r30']
HD[906] = 32'b001100_00001_10010_0000000000000000; //['load', '$r1', '$r18']
HD[907] = 32'b001101_10011_000000000000000000000; //['loadi', '$r19', '0']
HD[908] = 32'b011011_10100_00001_10011_00000000000; //['eq', '$r20', '$r1', '$r19']
HD[909] = 32'b100010_00000_10100_0000001110010001; //['jei', '$r0', '$r20', 'L29']
HD[910] = 32'b001101_11110_000000000000000001111; //['loadi', '$r30', 15]
HD[911] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[912] = 32'b001100_11011_00001_0000000000000000; //['load', '$r27', '$r1']
HD[913] = 32'b001101_11110_000000000000000010011; //['loadi', '$r30', 19]
HD[914] = 32'b000001_10011_11000_11110_00000000000; //['add', '$r19', '$r24', '$r30']
HD[915] = 32'b001100_00001_10011_0000000000000000; //['load', '$r1', '$r19']
HD[916] = 32'b001101_10100_000000000000000000001; //['loadi', '$r20', '1']
HD[917] = 32'b011011_10101_00001_10100_00000000000; //['eq', '$r21', '$r1', '$r20']
HD[918] = 32'b100010_00000_10101_0000001110011010; //['jei', '$r0', '$r21', 'L31']
HD[919] = 32'b001101_11110_000000000000000010000; //['loadi', '$r30', 16]
HD[920] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[921] = 32'b001100_11011_00001_0000000000000000; //['load', '$r27', '$r1']
HD[922] = 32'b001101_11110_000000000000000010011; //['loadi', '$r30', 19]
HD[923] = 32'b000001_10100_11000_11110_00000000000; //['add', '$r20', '$r24', '$r30']
HD[924] = 32'b001100_00001_10100_0000000000000000; //['load', '$r1', '$r20']
HD[925] = 32'b001101_10101_000000000000000000010; //['loadi', '$r21', '2']
HD[926] = 32'b011011_00001_00001_10101_00000000000; //['eq', '$r1', '$r1', '$r21']
HD[927] = 32'b100010_00000_00001_0000001110100011; //['jei', '$r0', '$r1', 'L33']
HD[928] = 32'b001101_11110_000000000000000010001; //['loadi', '$r30', 17]
HD[929] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[930] = 32'b001100_11011_00001_0000000000000000; //['load', '$r27', '$r1']
HD[931] = 32'b001101_11110_000000000000000010011; //['loadi', '$r30', 19]
HD[932] = 32'b000001_00010_11000_11110_00000000000; //['add', '$r2', '$r24', '$r30']
HD[933] = 32'b001100_00001_00010_0000000000000000; //['load', '$r1', '$r2']
HD[934] = 32'b001101_00011_000000000000000000011; //['loadi', '$r3', '3']
HD[935] = 32'b011011_00100_00001_00011_00000000000; //['eq', '$r4', '$r1', '$r3']
HD[936] = 32'b100010_00000_00100_0000001110101100; //['jei', '$r0', '$r4', 'L35']
HD[937] = 32'b001101_11110_000000000000000010010; //['loadi', '$r30', 18]
HD[938] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[939] = 32'b001100_11011_00001_0000000000000000; //['load', '$r27', '$r1']
HD[940] = 32'b101101_11011_000000000000000000000; //['setpcprog', '$r27']
HD[941] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[942] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[943] = 32'b011000_00000000000000000000000000; //['nop', ' ']
HD[944] = 32'b101011_00000000000000000000000000; //['setprogos', ' ']
HD[945] = 32'b011000_00000000000000000000000000; //['nop', ' ']
HD[946] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[947] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[948] = 32'b101100_00000000000000000000000000; //['savepcprog', ' ']
HD[949] = 32'b001101_11110_000000000000000010011; //['loadi', '$r30', 19]
HD[950] = 32'b000001_00011_11000_11110_00000000000; //['add', '$r3', '$r24', '$r30']
HD[951] = 32'b001100_00001_00011_0000000000000000; //['load', '$r1', '$r3']
HD[952] = 32'b001101_00100_000000000000000000000; //['loadi', '$r4', '0']
HD[953] = 32'b011011_00101_00001_00100_00000000000; //['eq', '$r5', '$r1', '$r4']
HD[954] = 32'b100010_00000_00101_0000001110111110; //['jei', '$r0', '$r5', 'L37']
HD[955] = 32'b001101_11110_000000000000000001111; //['loadi', '$r30', 15]
HD[956] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[957] = 32'b001110_11011_00001_0000000000000000; //['store', '$r27', '$r1']
HD[958] = 32'b001101_11110_000000000000000010011; //['loadi', '$r30', 19]
HD[959] = 32'b000001_00100_11000_11110_00000000000; //['add', '$r4', '$r24', '$r30']
HD[960] = 32'b001100_00001_00100_0000000000000000; //['load', '$r1', '$r4']
HD[961] = 32'b001101_00101_000000000000000000001; //['loadi', '$r5', '1']
HD[962] = 32'b011011_00110_00001_00101_00000000000; //['eq', '$r6', '$r1', '$r5']
HD[963] = 32'b100010_00000_00110_0000001111000111; //['jei', '$r0', '$r6', 'L39']
HD[964] = 32'b001101_11110_000000000000000010000; //['loadi', '$r30', 16]
HD[965] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[966] = 32'b001110_11011_00001_0000000000000000; //['store', '$r27', '$r1']
HD[967] = 32'b001101_11110_000000000000000010011; //['loadi', '$r30', 19]
HD[968] = 32'b000001_00101_11000_11110_00000000000; //['add', '$r5', '$r24', '$r30']
HD[969] = 32'b001100_00001_00101_0000000000000000; //['load', '$r1', '$r5']
HD[970] = 32'b001101_00110_000000000000000000010; //['loadi', '$r6', '2']
HD[971] = 32'b011011_00111_00001_00110_00000000000; //['eq', '$r7', '$r1', '$r6']
HD[972] = 32'b100010_00000_00111_0000001111010000; //['jei', '$r0', '$r7', 'L41']
HD[973] = 32'b001101_11110_000000000000000010001; //['loadi', '$r30', 17]
HD[974] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[975] = 32'b001110_11011_00001_0000000000000000; //['store', '$r27', '$r1']
HD[976] = 32'b001101_11110_000000000000000010011; //['loadi', '$r30', 19]
HD[977] = 32'b000001_00110_11000_11110_00000000000; //['add', '$r6', '$r24', '$r30']
HD[978] = 32'b001100_00001_00110_0000000000000000; //['load', '$r1', '$r6']
HD[979] = 32'b001101_00111_000000000000000000011; //['loadi', '$r7', '3']
HD[980] = 32'b011011_01000_00001_00111_00000000000; //['eq', '$r8', '$r1', '$r7']
HD[981] = 32'b100010_00000_01000_0000001111011001; //['jei', '$r0', '$r8', 'L43']
HD[982] = 32'b001101_11110_000000000000000010010; //['loadi', '$r30', 18]
HD[983] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[984] = 32'b001110_11011_00001_0000000000000000; //['store', '$r27', '$r1']
HD[985] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[986] = 32'b001111_11010_11010_0000000000000000; //['move', '$r26', '$r26']
HD[987] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[988] = 32'b001101_11110_000000000000000001010; //['loadi', '$r30', 10]
HD[989] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[990] = 32'b001110_11010_00001_0000000000000000; //['store', '$r26', '$r1']
HD[991] = 32'b001101_11110_000000000000000001010; //['loadi', '$r30', 10]
HD[992] = 32'b000001_00111_11000_11110_00000000000; //['add', '$r7', '$r24', '$r30']
HD[993] = 32'b001100_00001_00111_0000000000000000; //['load', '$r1', '$r7']
HD[994] = 32'b010111_00001_000000000000000000000; //['out', '$r1']
HD[995] = 32'b001101_11110_000000000000000001010; //['loadi', '$r30', 10]
HD[996] = 32'b000001_00111_11000_11110_00000000000; //['add', '$r7', '$r24', '$r30']
HD[997] = 32'b001100_00001_00111_0000000000000000; //['load', '$r1', '$r7']
HD[998] = 32'b001101_01000_000000000000000000000; //['loadi', '$r8', '0']
HD[999] = 32'b011011_01001_00001_01000_00000000000; //['eq', '$r9', '$r1', '$r8']
HD[1000] = 32'b100010_00000_01001_0000001111110001; //['jei', '$r0', '$r9', 'L45']
HD[1001] = 32'b001101_01000_000000000000000000000; //['loadi', '$r8', 0]
HD[1002] = 32'b000001_00001_11000_01000_00000000000; //['add', '$r1', '$r24', '$r8']
HD[1003] = 32'b001101_11110_000000000000000010011; //['loadi', '$r30', 19]
HD[1004] = 32'b000001_01000_11000_11110_00000000000; //['add', '$r8', '$r24', '$r30']
HD[1005] = 32'b001100_01001_01000_0000000000000000; //['load', '$r9', '$r8']
HD[1006] = 32'b000001_10101_00001_01001_00000000000; //['add', '$r21', '$r1', '$r9']
HD[1007] = 32'b001101_00001_000000000000000000000; //['loadi', '$r1', '0']
HD[1008] = 32'b001110_00001_10101_0000000000000000; //['store', '$r1', '$r21']
HD[1009] = 32'b001101_11110_000000000000000001010; //['loadi', '$r30', 10]
HD[1010] = 32'b000001_01000_11000_11110_00000000000; //['add', '$r8', '$r24', '$r30']
HD[1011] = 32'b001100_00001_01000_0000000000000000; //['load', '$r1', '$r8']
HD[1012] = 32'b001101_01001_000000000000000000001; //['loadi', '$r9', '1']
HD[1013] = 32'b011011_10101_00001_01001_00000000000; //['eq', '$r21', '$r1', '$r9']
HD[1014] = 32'b100010_00000_10101_0000010000001111; //['jei', '$r0', '$r21', 'L47']
HD[1015] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1016] = 32'b001111_11001_11001_0000000000000000; //['move', '$r25', '$r25']
HD[1017] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1018] = 32'b001101_11110_000000000000000001011; //['loadi', '$r30', 11]
HD[1019] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[1020] = 32'b001110_11001_00001_0000000000000000; //['store', '$r25', '$r1']
HD[1021] = 32'b001101_11110_000000000000000010011; //['loadi', '$r30', 19]
HD[1022] = 32'b000001_01001_11000_11110_00000000000; //['add', '$r9', '$r24', '$r30']
HD[1023] = 32'b001100_00001_01001_0000000000000000; //['load', '$r1', '$r9']
HD[1024] = 32'b010111_00001_000000000000000000000; //['out', '$r1']
HD[1025] = 32'b001101_11110_000000000000000001011; //['loadi', '$r30', 11]
HD[1026] = 32'b000001_01001_11000_11110_00000000000; //['add', '$r9', '$r24', '$r30']
HD[1027] = 32'b001100_00001_01001_0000000000000000; //['load', '$r1', '$r9']
HD[1028] = 32'b010111_00001_000000000000000000000; //['out', '$r1']
HD[1029] = 32'b001101_11110_000000000000000001010; //['loadi', '$r30', 10]
HD[1030] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[1031] = 32'b001101_10101_000000000000000000000; //['loadi', '$r21', '0']
HD[1032] = 32'b001110_10101_00001_0000000000000000; //['store', '$r21', '$r1']
HD[1033] = 32'b001101_11110_000000000000000001010; //['loadi', '$r30', 10]
HD[1034] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[1035] = 32'b001100_11010_00001_0000000000000000; //['load', '$r26', '$r1']
HD[1036] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[1037] = 32'b001111_11010_11010_0000000000000000; //['move', '$r26', '$r26']
HD[1038] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[1039] = 32'b001101_11110_000000000000000001010; //['loadi', '$r30', 10]
HD[1040] = 32'b000001_01001_11000_11110_00000000000; //['add', '$r9', '$r24', '$r30']
HD[1041] = 32'b001100_00001_01001_0000000000000000; //['load', '$r1', '$r9']
HD[1042] = 32'b001101_10101_000000000000000000010; //['loadi', '$r21', '2']
HD[1043] = 32'b011011_00001_00001_10101_00000000000; //['eq', '$r1', '$r1', '$r21']
HD[1044] = 32'b100010_00000_00001_0000010000101110; //['jei', '$r0', '$r1', 'L49']
HD[1045] = 32'b001101_11110_000000000000000010011; //['loadi', '$r30', 19]
HD[1046] = 32'b000001_00010_11000_11110_00000000000; //['add', '$r2', '$r24', '$r30']
HD[1047] = 32'b001100_00001_00010_0000000000000000; //['load', '$r1', '$r2']
HD[1048] = 32'b010111_00001_000000000000000000000; //['out', '$r1']
HD[1049] = 32'b010110_11100_000000000000000000000; //['in', '$r28']
HD[1050] = 32'b001111_00001_11100_0000000000000000; //['move', '$r1', '$r28']
HD[1051] = 32'b001101_11110_000000000000000001100; //['loadi', '$r30', 12]
HD[1052] = 32'b000001_00010_11000_11110_00000000000; //['add', '$r2', '$r24', '$r30']
HD[1053] = 32'b001110_00001_00010_0000000000000000; //['store', '$r1', '$r2']
HD[1054] = 32'b001101_11110_000000000000000001100; //['loadi', '$r30', 12]
HD[1055] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[1056] = 32'b001100_11100_00001_0000000000000000; //['load', '$r28', '$r1']
HD[1057] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[1058] = 32'b001111_11100_11100_0000000000000000; //['move', '$r28', '$r28']
HD[1059] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[1060] = 32'b001101_11110_000000000000000001010; //['loadi', '$r30', 10]
HD[1061] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[1062] = 32'b001101_00011_000000000000000000000; //['loadi', '$r3', '0']
HD[1063] = 32'b001110_00011_00001_0000000000000000; //['store', '$r3', '$r1']
HD[1064] = 32'b001101_11110_000000000000000001010; //['loadi', '$r30', 10]
HD[1065] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[1066] = 32'b001100_11010_00001_0000000000000000; //['load', '$r26', '$r1']
HD[1067] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[1068] = 32'b001111_11010_11010_0000000000000000; //['move', '$r26', '$r26']
HD[1069] = 32'b100101_00000000000000000000000000; //['flagrd', ' ']
HD[1070] = 32'b001101_11110_000000000000000010011; //['loadi', '$r30', 19]
HD[1071] = 32'b000001_00010_11000_11110_00000000000; //['add', '$r2', '$r24', '$r30']
HD[1072] = 32'b001100_00001_00010_0000000000000000; //['load', '$r1', '$r2']
HD[1073] = 32'b001101_00011_000000000000000000000; //['loadi', '$r3', '0']
HD[1074] = 32'b011011_00100_00001_00011_00000000000; //['eq', '$r4', '$r1', '$r3']
HD[1075] = 32'b100010_00000_00100_0000010011010100; //['jei', '$r0', '$r4', 'L51']
HD[1076] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1077] = 32'b001111_10110_00000_0000000000000000; //['move', '$r22', '$r0']
HD[1078] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1079] = 32'b001101_00001_000000000000110010000; //['loadi', '$r1', '400']
HD[1080] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1081] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1082] = 32'b001111_10110_00001_0000000000000000; //['move', '$r22', '$r1']
HD[1083] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1084] = 32'b001101_00001_000000000000110010001; //['loadi', '$r1', '401']
HD[1085] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1086] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1087] = 32'b001111_10110_00010_0000000000000000; //['move', '$r22', '$r2']
HD[1088] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1089] = 32'b001101_00001_000000000000110010010; //['loadi', '$r1', '402']
HD[1090] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1091] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1092] = 32'b001111_10110_00011_0000000000000000; //['move', '$r22', '$r3']
HD[1093] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1094] = 32'b001101_00001_000000000000110010011; //['loadi', '$r1', '403']
HD[1095] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1096] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1097] = 32'b001111_10110_00100_0000000000000000; //['move', '$r22', '$r4']
HD[1098] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1099] = 32'b001101_00001_000000000000110010100; //['loadi', '$r1', '404']
HD[1100] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1101] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1102] = 32'b001111_10110_00101_0000000000000000; //['move', '$r22', '$r5']
HD[1103] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1104] = 32'b001101_00001_000000000000110010101; //['loadi', '$r1', '405']
HD[1105] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1106] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1107] = 32'b001111_10110_00110_0000000000000000; //['move', '$r22', '$r6']
HD[1108] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1109] = 32'b001101_00001_000000000000110010110; //['loadi', '$r1', '406']
HD[1110] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1111] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1112] = 32'b001111_10110_00111_0000000000000000; //['move', '$r22', '$r7']
HD[1113] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1114] = 32'b001101_00001_000000000000110010111; //['loadi', '$r1', '407']
HD[1115] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1116] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1117] = 32'b001111_10110_01000_0000000000000000; //['move', '$r22', '$r8']
HD[1118] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1119] = 32'b001101_00001_000000000000110011000; //['loadi', '$r1', '408']
HD[1120] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1121] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1122] = 32'b001111_10110_01001_0000000000000000; //['move', '$r22', '$r9']
HD[1123] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1124] = 32'b001101_00001_000000000000110011001; //['loadi', '$r1', '409']
HD[1125] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1126] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1127] = 32'b001111_10110_01010_0000000000000000; //['move', '$r22', '$r10']
HD[1128] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1129] = 32'b001101_00001_000000000000110011010; //['loadi', '$r1', '410']
HD[1130] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1131] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1132] = 32'b001111_10110_01011_0000000000000000; //['move', '$r22', '$r11']
HD[1133] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1134] = 32'b001101_00001_000000000000110011011; //['loadi', '$r1', '411']
HD[1135] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1136] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1137] = 32'b001111_10110_01100_0000000000000000; //['move', '$r22', '$r12']
HD[1138] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1139] = 32'b001101_00001_000000000000110011100; //['loadi', '$r1', '412']
HD[1140] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1141] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1142] = 32'b001111_10110_01101_0000000000000000; //['move', '$r22', '$r13']
HD[1143] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1144] = 32'b001101_00001_000000000000110011101; //['loadi', '$r1', '413']
HD[1145] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1146] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1147] = 32'b001111_10110_01110_0000000000000000; //['move', '$r22', '$r14']
HD[1148] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1149] = 32'b001101_00001_000000000000110011110; //['loadi', '$r1', '414']
HD[1150] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1151] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1152] = 32'b001111_10110_01111_0000000000000000; //['move', '$r22', '$r15']
HD[1153] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1154] = 32'b001101_00001_000000000000110011111; //['loadi', '$r1', '415']
HD[1155] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1156] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1157] = 32'b001111_10110_10000_0000000000000000; //['move', '$r22', '$r16']
HD[1158] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1159] = 32'b001101_00001_000000000000110100000; //['loadi', '$r1', '416']
HD[1160] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1161] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1162] = 32'b001111_10110_10001_0000000000000000; //['move', '$r22', '$r17']
HD[1163] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1164] = 32'b001101_00001_000000000000110100001; //['loadi', '$r1', '417']
HD[1165] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1166] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1167] = 32'b001111_10110_10010_0000000000000000; //['move', '$r22', '$r18']
HD[1168] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1169] = 32'b001101_00001_000000000000110100010; //['loadi', '$r1', '418']
HD[1170] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1171] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1172] = 32'b001111_10110_10011_0000000000000000; //['move', '$r22', '$r19']
HD[1173] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1174] = 32'b001101_00001_000000000000110100011; //['loadi', '$r1', '419']
HD[1175] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1176] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1177] = 32'b001111_10110_10100_0000000000000000; //['move', '$r22', '$r20']
HD[1178] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1179] = 32'b001101_00001_000000000000110100100; //['loadi', '$r1', '420']
HD[1180] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1181] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1182] = 32'b001111_10110_10101_0000000000000000; //['move', '$r22', '$r21']
HD[1183] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1184] = 32'b001101_00001_000000000000110100101; //['loadi', '$r1', '421']
HD[1185] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1186] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1187] = 32'b001111_10110_10110_0000000000000000; //['move', '$r22', '$r22']
HD[1188] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1189] = 32'b001101_00001_000000000000110100110; //['loadi', '$r1', '422']
HD[1190] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1191] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1192] = 32'b001111_10110_10111_0000000000000000; //['move', '$r22', '$r23']
HD[1193] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1194] = 32'b001101_00001_000000000000110100111; //['loadi', '$r1', '423']
HD[1195] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1196] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1197] = 32'b001111_10110_11000_0000000000000000; //['move', '$r22', '$r24']
HD[1198] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1199] = 32'b001101_00001_000000000000110101000; //['loadi', '$r1', '424']
HD[1200] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1201] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1202] = 32'b001111_10110_11001_0000000000000000; //['move', '$r22', '$r25']
HD[1203] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1204] = 32'b001101_00001_000000000000110101001; //['loadi', '$r1', '425']
HD[1205] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1206] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1207] = 32'b001111_10110_11010_0000000000000000; //['move', '$r22', '$r26']
HD[1208] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1209] = 32'b001101_00001_000000000000110101010; //['loadi', '$r1', '426']
HD[1210] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1211] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1212] = 32'b001111_10110_11011_0000000000000000; //['move', '$r22', '$r27']
HD[1213] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1214] = 32'b001101_00001_000000000000110101011; //['loadi', '$r1', '427']
HD[1215] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1216] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1217] = 32'b001111_10110_11100_0000000000000000; //['move', '$r22', '$r28']
HD[1218] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1219] = 32'b001101_00001_000000000000110101100; //['loadi', '$r1', '428']
HD[1220] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1221] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1222] = 32'b001111_10110_11101_0000000000000000; //['move', '$r22', '$r29']
HD[1223] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1224] = 32'b001101_00001_000000000000110101101; //['loadi', '$r1', '429']
HD[1225] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1226] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1227] = 32'b001111_10110_11110_0000000000000000; //['move', '$r22', '$r30']
HD[1228] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1229] = 32'b001101_00001_000000000000110101110; //['loadi', '$r1', '430']
HD[1230] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1231] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1232] = 32'b001111_10110_11111_0000000000000000; //['move', '$r22', '$r31']
HD[1233] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1234] = 32'b001101_00001_000000000000110101111; //['loadi', '$r1', '431']
HD[1235] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1236] = 32'b001101_11110_000000000000000010011; //['loadi', '$r30', 19]
HD[1237] = 32'b000001_00011_11000_11110_00000000000; //['add', '$r3', '$r24', '$r30']
HD[1238] = 32'b001100_00001_00011_0000000000000000; //['load', '$r1', '$r3']
HD[1239] = 32'b001101_00100_000000000000000000001; //['loadi', '$r4', '1']
HD[1240] = 32'b011011_00101_00001_00100_00000000000; //['eq', '$r5', '$r1', '$r4']
HD[1241] = 32'b100010_00000_00101_0000010101111010; //['jei', '$r0', '$r5', 'L53']
HD[1242] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1243] = 32'b001111_10110_00000_0000000000000000; //['move', '$r22', '$r0']
HD[1244] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1245] = 32'b001101_00001_000000000000110110000; //['loadi', '$r1', '432']
HD[1246] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1247] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1248] = 32'b001111_10110_00001_0000000000000000; //['move', '$r22', '$r1']
HD[1249] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1250] = 32'b001101_00001_000000000000110110001; //['loadi', '$r1', '433']
HD[1251] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1252] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1253] = 32'b001111_10110_00010_0000000000000000; //['move', '$r22', '$r2']
HD[1254] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1255] = 32'b001101_00001_000000000000110110010; //['loadi', '$r1', '434']
HD[1256] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1257] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1258] = 32'b001111_10110_00011_0000000000000000; //['move', '$r22', '$r3']
HD[1259] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1260] = 32'b001101_00001_000000000000110110011; //['loadi', '$r1', '435']
HD[1261] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1262] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1263] = 32'b001111_10110_00100_0000000000000000; //['move', '$r22', '$r4']
HD[1264] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1265] = 32'b001101_00001_000000000000110110100; //['loadi', '$r1', '436']
HD[1266] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1267] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1268] = 32'b001111_10110_00101_0000000000000000; //['move', '$r22', '$r5']
HD[1269] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1270] = 32'b001101_00001_000000000000110110101; //['loadi', '$r1', '437']
HD[1271] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1272] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1273] = 32'b001111_10110_00110_0000000000000000; //['move', '$r22', '$r6']
HD[1274] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1275] = 32'b001101_00001_000000000000110110110; //['loadi', '$r1', '438']
HD[1276] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1277] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1278] = 32'b001111_10110_00111_0000000000000000; //['move', '$r22', '$r7']
HD[1279] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1280] = 32'b001101_00001_000000000000110110111; //['loadi', '$r1', '439']
HD[1281] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1282] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1283] = 32'b001111_10110_01000_0000000000000000; //['move', '$r22', '$r8']
HD[1284] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1285] = 32'b001101_00001_000000000000110111000; //['loadi', '$r1', '440']
HD[1286] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1287] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1288] = 32'b001111_10110_01001_0000000000000000; //['move', '$r22', '$r9']
HD[1289] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1290] = 32'b001101_00001_000000000000110111001; //['loadi', '$r1', '441']
HD[1291] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1292] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1293] = 32'b001111_10110_01010_0000000000000000; //['move', '$r22', '$r10']
HD[1294] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1295] = 32'b001101_00001_000000000000110111010; //['loadi', '$r1', '442']
HD[1296] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1297] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1298] = 32'b001111_10110_01011_0000000000000000; //['move', '$r22', '$r11']
HD[1299] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1300] = 32'b001101_00001_000000000000110111011; //['loadi', '$r1', '443']
HD[1301] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1302] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1303] = 32'b001111_10110_01100_0000000000000000; //['move', '$r22', '$r12']
HD[1304] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1305] = 32'b001101_00001_000000000000110111100; //['loadi', '$r1', '444']
HD[1306] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1307] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1308] = 32'b001111_10110_01101_0000000000000000; //['move', '$r22', '$r13']
HD[1309] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1310] = 32'b001101_00001_000000000000110111101; //['loadi', '$r1', '445']
HD[1311] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1312] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1313] = 32'b001111_10110_01110_0000000000000000; //['move', '$r22', '$r14']
HD[1314] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1315] = 32'b001101_00001_000000000000110111110; //['loadi', '$r1', '446']
HD[1316] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1317] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1318] = 32'b001111_10110_01111_0000000000000000; //['move', '$r22', '$r15']
HD[1319] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1320] = 32'b001101_00001_000000000000110111111; //['loadi', '$r1', '447']
HD[1321] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1322] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1323] = 32'b001111_10110_10000_0000000000000000; //['move', '$r22', '$r16']
HD[1324] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1325] = 32'b001101_00001_000000000000111000000; //['loadi', '$r1', '448']
HD[1326] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1327] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1328] = 32'b001111_10110_10001_0000000000000000; //['move', '$r22', '$r17']
HD[1329] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1330] = 32'b001101_00001_000000000000111000001; //['loadi', '$r1', '449']
HD[1331] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1332] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1333] = 32'b001111_10110_10010_0000000000000000; //['move', '$r22', '$r18']
HD[1334] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1335] = 32'b001101_00001_000000000000111000010; //['loadi', '$r1', '450']
HD[1336] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1337] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1338] = 32'b001111_10110_10011_0000000000000000; //['move', '$r22', '$r19']
HD[1339] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1340] = 32'b001101_00001_000000000000111000011; //['loadi', '$r1', '451']
HD[1341] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1342] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1343] = 32'b001111_10110_10100_0000000000000000; //['move', '$r22', '$r20']
HD[1344] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1345] = 32'b001101_00001_000000000000111000100; //['loadi', '$r1', '452']
HD[1346] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1347] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1348] = 32'b001111_10110_10101_0000000000000000; //['move', '$r22', '$r21']
HD[1349] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1350] = 32'b001101_00001_000000000000111000101; //['loadi', '$r1', '453']
HD[1351] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1352] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1353] = 32'b001111_10110_10110_0000000000000000; //['move', '$r22', '$r22']
HD[1354] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1355] = 32'b001101_00001_000000000000111000110; //['loadi', '$r1', '454']
HD[1356] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1357] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1358] = 32'b001111_10110_10111_0000000000000000; //['move', '$r22', '$r23']
HD[1359] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1360] = 32'b001101_00001_000000000000111000111; //['loadi', '$r1', '455']
HD[1361] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1362] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1363] = 32'b001111_10110_11000_0000000000000000; //['move', '$r22', '$r24']
HD[1364] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1365] = 32'b001101_00001_000000000000111001000; //['loadi', '$r1', '456']
HD[1366] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1367] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1368] = 32'b001111_10110_11001_0000000000000000; //['move', '$r22', '$r25']
HD[1369] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1370] = 32'b001101_00001_000000000000111001001; //['loadi', '$r1', '457']
HD[1371] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1372] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1373] = 32'b001111_10110_11010_0000000000000000; //['move', '$r22', '$r26']
HD[1374] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1375] = 32'b001101_00001_000000000000111001010; //['loadi', '$r1', '458']
HD[1376] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1377] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1378] = 32'b001111_10110_11011_0000000000000000; //['move', '$r22', '$r27']
HD[1379] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1380] = 32'b001101_00001_000000000000111001011; //['loadi', '$r1', '459']
HD[1381] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1382] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1383] = 32'b001111_10110_11100_0000000000000000; //['move', '$r22', '$r28']
HD[1384] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1385] = 32'b001101_00001_000000000000111001100; //['loadi', '$r1', '460']
HD[1386] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1387] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1388] = 32'b001111_10110_11101_0000000000000000; //['move', '$r22', '$r29']
HD[1389] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1390] = 32'b001101_00001_000000000000111001101; //['loadi', '$r1', '461']
HD[1391] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1392] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1393] = 32'b001111_10110_11110_0000000000000000; //['move', '$r22', '$r30']
HD[1394] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1395] = 32'b001101_00001_000000000000111001110; //['loadi', '$r1', '462']
HD[1396] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1397] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1398] = 32'b001111_10110_11111_0000000000000000; //['move', '$r22', '$r31']
HD[1399] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1400] = 32'b001101_00001_000000000000111001111; //['loadi', '$r1', '463']
HD[1401] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1402] = 32'b001101_11110_000000000000000010011; //['loadi', '$r30', 19]
HD[1403] = 32'b000001_00100_11000_11110_00000000000; //['add', '$r4', '$r24', '$r30']
HD[1404] = 32'b001100_00001_00100_0000000000000000; //['load', '$r1', '$r4']
HD[1405] = 32'b001101_00101_000000000000000000010; //['loadi', '$r5', '2']
HD[1406] = 32'b011011_00110_00001_00101_00000000000; //['eq', '$r6', '$r1', '$r5']
HD[1407] = 32'b100010_00000_00110_0000011000100000; //['jei', '$r0', '$r6', 'L55']
HD[1408] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1409] = 32'b001111_10110_00000_0000000000000000; //['move', '$r22', '$r0']
HD[1410] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1411] = 32'b001101_00001_000000000000100101100; //['loadi', '$r1', '300']
HD[1412] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1413] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1414] = 32'b001111_10110_00001_0000000000000000; //['move', '$r22', '$r1']
HD[1415] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1416] = 32'b001101_00001_000000000000100101101; //['loadi', '$r1', '301']
HD[1417] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1418] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1419] = 32'b001111_10110_00010_0000000000000000; //['move', '$r22', '$r2']
HD[1420] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1421] = 32'b001101_00001_000000000000100101110; //['loadi', '$r1', '302']
HD[1422] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1423] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1424] = 32'b001111_10110_00011_0000000000000000; //['move', '$r22', '$r3']
HD[1425] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1426] = 32'b001101_00001_000000000000100101111; //['loadi', '$r1', '303']
HD[1427] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1428] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1429] = 32'b001111_10110_00100_0000000000000000; //['move', '$r22', '$r4']
HD[1430] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1431] = 32'b001101_00001_000000000000100110000; //['loadi', '$r1', '304']
HD[1432] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1433] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1434] = 32'b001111_10110_00101_0000000000000000; //['move', '$r22', '$r5']
HD[1435] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1436] = 32'b001101_00001_000000000000100110001; //['loadi', '$r1', '305']
HD[1437] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1438] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1439] = 32'b001111_10110_00110_0000000000000000; //['move', '$r22', '$r6']
HD[1440] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1441] = 32'b001101_00001_000000000000100110010; //['loadi', '$r1', '306']
HD[1442] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1443] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1444] = 32'b001111_10110_00111_0000000000000000; //['move', '$r22', '$r7']
HD[1445] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1446] = 32'b001101_00001_000000000000100110011; //['loadi', '$r1', '307']
HD[1447] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1448] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1449] = 32'b001111_10110_01000_0000000000000000; //['move', '$r22', '$r8']
HD[1450] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1451] = 32'b001101_00001_000000000000100110100; //['loadi', '$r1', '308']
HD[1452] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1453] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1454] = 32'b001111_10110_01001_0000000000000000; //['move', '$r22', '$r9']
HD[1455] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1456] = 32'b001101_00001_000000000000100110101; //['loadi', '$r1', '309']
HD[1457] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1458] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1459] = 32'b001111_10110_01010_0000000000000000; //['move', '$r22', '$r10']
HD[1460] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1461] = 32'b001101_00001_000000000000100110110; //['loadi', '$r1', '310']
HD[1462] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1463] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1464] = 32'b001111_10110_01011_0000000000000000; //['move', '$r22', '$r11']
HD[1465] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1466] = 32'b001101_00001_000000000000100110111; //['loadi', '$r1', '311']
HD[1467] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1468] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1469] = 32'b001111_10110_01100_0000000000000000; //['move', '$r22', '$r12']
HD[1470] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1471] = 32'b001101_00001_000000000000100111000; //['loadi', '$r1', '312']
HD[1472] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1473] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1474] = 32'b001111_10110_01101_0000000000000000; //['move', '$r22', '$r13']
HD[1475] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1476] = 32'b001101_00001_000000000000100111001; //['loadi', '$r1', '313']
HD[1477] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1478] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1479] = 32'b001111_10110_01110_0000000000000000; //['move', '$r22', '$r14']
HD[1480] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1481] = 32'b001101_00001_000000000000100111010; //['loadi', '$r1', '314']
HD[1482] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1483] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1484] = 32'b001111_10110_01111_0000000000000000; //['move', '$r22', '$r15']
HD[1485] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1486] = 32'b001101_00001_000000000000100111011; //['loadi', '$r1', '315']
HD[1487] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1488] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1489] = 32'b001111_10110_10000_0000000000000000; //['move', '$r22', '$r16']
HD[1490] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1491] = 32'b001101_00001_000000000000100111100; //['loadi', '$r1', '316']
HD[1492] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1493] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1494] = 32'b001111_10110_10001_0000000000000000; //['move', '$r22', '$r17']
HD[1495] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1496] = 32'b001101_00001_000000000000100111101; //['loadi', '$r1', '317']
HD[1497] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1498] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1499] = 32'b001111_10110_10010_0000000000000000; //['move', '$r22', '$r18']
HD[1500] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1501] = 32'b001101_00001_000000000000100111110; //['loadi', '$r1', '318']
HD[1502] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1503] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1504] = 32'b001111_10110_10011_0000000000000000; //['move', '$r22', '$r19']
HD[1505] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1506] = 32'b001101_00001_000000000000100111111; //['loadi', '$r1', '319']
HD[1507] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1508] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1509] = 32'b001111_10110_10100_0000000000000000; //['move', '$r22', '$r20']
HD[1510] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1511] = 32'b001101_00001_000000000000101000000; //['loadi', '$r1', '320']
HD[1512] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1513] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1514] = 32'b001111_10110_10101_0000000000000000; //['move', '$r22', '$r21']
HD[1515] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1516] = 32'b001101_00001_000000000000101000001; //['loadi', '$r1', '321']
HD[1517] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1518] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1519] = 32'b001111_10110_10110_0000000000000000; //['move', '$r22', '$r22']
HD[1520] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1521] = 32'b001101_00001_000000000000101000010; //['loadi', '$r1', '322']
HD[1522] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1523] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1524] = 32'b001111_10110_10111_0000000000000000; //['move', '$r22', '$r23']
HD[1525] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1526] = 32'b001101_00001_000000000000101000011; //['loadi', '$r1', '323']
HD[1527] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1528] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1529] = 32'b001111_10110_11000_0000000000000000; //['move', '$r22', '$r24']
HD[1530] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1531] = 32'b001101_00001_000000000000101000100; //['loadi', '$r1', '324']
HD[1532] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1533] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1534] = 32'b001111_10110_11001_0000000000000000; //['move', '$r22', '$r25']
HD[1535] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1536] = 32'b001101_00001_000000000000101000101; //['loadi', '$r1', '325']
HD[1537] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1538] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1539] = 32'b001111_10110_11010_0000000000000000; //['move', '$r22', '$r26']
HD[1540] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1541] = 32'b001101_00001_000000000000101000110; //['loadi', '$r1', '326']
HD[1542] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1543] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1544] = 32'b001111_10110_11011_0000000000000000; //['move', '$r22', '$r27']
HD[1545] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1546] = 32'b001101_00001_000000000000101000111; //['loadi', '$r1', '327']
HD[1547] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1548] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1549] = 32'b001111_10110_11100_0000000000000000; //['move', '$r22', '$r28']
HD[1550] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1551] = 32'b001101_00001_000000000000101001000; //['loadi', '$r1', '328']
HD[1552] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1553] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1554] = 32'b001111_10110_11101_0000000000000000; //['move', '$r22', '$r29']
HD[1555] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1556] = 32'b001101_00001_000000000000101001001; //['loadi', '$r1', '329']
HD[1557] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1558] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1559] = 32'b001111_10110_11110_0000000000000000; //['move', '$r22', '$r30']
HD[1560] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1561] = 32'b001101_00001_000000000000101001010; //['loadi', '$r1', '330']
HD[1562] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1563] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1564] = 32'b001111_10110_11111_0000000000000000; //['move', '$r22', '$r31']
HD[1565] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1566] = 32'b001101_00001_000000000000101001011; //['loadi', '$r1', '331']
HD[1567] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1568] = 32'b001101_11110_000000000000000010011; //['loadi', '$r30', 19]
HD[1569] = 32'b000001_00101_11000_11110_00000000000; //['add', '$r5', '$r24', '$r30']
HD[1570] = 32'b001100_00001_00101_0000000000000000; //['load', '$r1', '$r5']
HD[1571] = 32'b001101_00110_000000000000000000011; //['loadi', '$r6', '3']
HD[1572] = 32'b011011_00111_00001_00110_00000000000; //['eq', '$r7', '$r1', '$r6']
HD[1573] = 32'b100010_00000_00111_0000011011000110; //['jei', '$r0', '$r7', 'L57']
HD[1574] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1575] = 32'b001111_10110_00000_0000000000000000; //['move', '$r22', '$r0']
HD[1576] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1577] = 32'b001101_00001_000000000000101001100; //['loadi', '$r1', '332']
HD[1578] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1579] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1580] = 32'b001111_10110_00001_0000000000000000; //['move', '$r22', '$r1']
HD[1581] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1582] = 32'b001101_00001_000000000000101001101; //['loadi', '$r1', '333']
HD[1583] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1584] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1585] = 32'b001111_10110_00010_0000000000000000; //['move', '$r22', '$r2']
HD[1586] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1587] = 32'b001101_00001_000000000000101001110; //['loadi', '$r1', '334']
HD[1588] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1589] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1590] = 32'b001111_10110_00011_0000000000000000; //['move', '$r22', '$r3']
HD[1591] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1592] = 32'b001101_00001_000000000000101001111; //['loadi', '$r1', '335']
HD[1593] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1594] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1595] = 32'b001111_10110_00100_0000000000000000; //['move', '$r22', '$r4']
HD[1596] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1597] = 32'b001101_00001_000000000000101010000; //['loadi', '$r1', '336']
HD[1598] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1599] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1600] = 32'b001111_10110_00101_0000000000000000; //['move', '$r22', '$r5']
HD[1601] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1602] = 32'b001101_00001_000000000000101010001; //['loadi', '$r1', '337']
HD[1603] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1604] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1605] = 32'b001111_10110_00110_0000000000000000; //['move', '$r22', '$r6']
HD[1606] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1607] = 32'b001101_00001_000000000000101010010; //['loadi', '$r1', '338']
HD[1608] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1609] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1610] = 32'b001111_10110_00111_0000000000000000; //['move', '$r22', '$r7']
HD[1611] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1612] = 32'b001101_00001_000000000000101010011; //['loadi', '$r1', '339']
HD[1613] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1614] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1615] = 32'b001111_10110_01000_0000000000000000; //['move', '$r22', '$r8']
HD[1616] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1617] = 32'b001101_00001_000000000000101010100; //['loadi', '$r1', '340']
HD[1618] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1619] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1620] = 32'b001111_10110_01001_0000000000000000; //['move', '$r22', '$r9']
HD[1621] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1622] = 32'b001101_00001_000000000000101010101; //['loadi', '$r1', '341']
HD[1623] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1624] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1625] = 32'b001111_10110_01010_0000000000000000; //['move', '$r22', '$r10']
HD[1626] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1627] = 32'b001101_00001_000000000000101010110; //['loadi', '$r1', '342']
HD[1628] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1629] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1630] = 32'b001111_10110_01011_0000000000000000; //['move', '$r22', '$r11']
HD[1631] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1632] = 32'b001101_00001_000000000000101010111; //['loadi', '$r1', '343']
HD[1633] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1634] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1635] = 32'b001111_10110_01100_0000000000000000; //['move', '$r22', '$r12']
HD[1636] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1637] = 32'b001101_00001_000000000000101011000; //['loadi', '$r1', '344']
HD[1638] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1639] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1640] = 32'b001111_10110_01101_0000000000000000; //['move', '$r22', '$r13']
HD[1641] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1642] = 32'b001101_00001_000000000000101011001; //['loadi', '$r1', '345']
HD[1643] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1644] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1645] = 32'b001111_10110_01110_0000000000000000; //['move', '$r22', '$r14']
HD[1646] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1647] = 32'b001101_00001_000000000000101011010; //['loadi', '$r1', '346']
HD[1648] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1649] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1650] = 32'b001111_10110_01111_0000000000000000; //['move', '$r22', '$r15']
HD[1651] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1652] = 32'b001101_00001_000000000000101011011; //['loadi', '$r1', '347']
HD[1653] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1654] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1655] = 32'b001111_10110_10000_0000000000000000; //['move', '$r22', '$r16']
HD[1656] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1657] = 32'b001101_00001_000000000000101011100; //['loadi', '$r1', '348']
HD[1658] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1659] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1660] = 32'b001111_10110_10001_0000000000000000; //['move', '$r22', '$r17']
HD[1661] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1662] = 32'b001101_00001_000000000000101011101; //['loadi', '$r1', '349']
HD[1663] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1664] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1665] = 32'b001111_10110_10010_0000000000000000; //['move', '$r22', '$r18']
HD[1666] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1667] = 32'b001101_00001_000000000000101011110; //['loadi', '$r1', '350']
HD[1668] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1669] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1670] = 32'b001111_10110_10011_0000000000000000; //['move', '$r22', '$r19']
HD[1671] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1672] = 32'b001101_00001_000000000000101011111; //['loadi', '$r1', '351']
HD[1673] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1674] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1675] = 32'b001111_10110_10100_0000000000000000; //['move', '$r22', '$r20']
HD[1676] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1677] = 32'b001101_00001_000000000000101100000; //['loadi', '$r1', '352']
HD[1678] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1679] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1680] = 32'b001111_10110_10101_0000000000000000; //['move', '$r22', '$r21']
HD[1681] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1682] = 32'b001101_00001_000000000000101100001; //['loadi', '$r1', '353']
HD[1683] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1684] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1685] = 32'b001111_10110_10110_0000000000000000; //['move', '$r22', '$r22']
HD[1686] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1687] = 32'b001101_00001_000000000000101100010; //['loadi', '$r1', '354']
HD[1688] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1689] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1690] = 32'b001111_10110_10111_0000000000000000; //['move', '$r22', '$r23']
HD[1691] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1692] = 32'b001101_00001_000000000000101100011; //['loadi', '$r1', '355']
HD[1693] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1694] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1695] = 32'b001111_10110_11000_0000000000000000; //['move', '$r22', '$r24']
HD[1696] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1697] = 32'b001101_00001_000000000000101100100; //['loadi', '$r1', '356']
HD[1698] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1699] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1700] = 32'b001111_10110_11001_0000000000000000; //['move', '$r22', '$r25']
HD[1701] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1702] = 32'b001101_00001_000000000000101100101; //['loadi', '$r1', '357']
HD[1703] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1704] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1705] = 32'b001111_10110_11010_0000000000000000; //['move', '$r22', '$r26']
HD[1706] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1707] = 32'b001101_00001_000000000000101100110; //['loadi', '$r1', '358']
HD[1708] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1709] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1710] = 32'b001111_10110_11011_0000000000000000; //['move', '$r22', '$r27']
HD[1711] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1712] = 32'b001101_00001_000000000000101100111; //['loadi', '$r1', '359']
HD[1713] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1714] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1715] = 32'b001111_10110_11100_0000000000000000; //['move', '$r22', '$r28']
HD[1716] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1717] = 32'b001101_00001_000000000000101101000; //['loadi', '$r1', '360']
HD[1718] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1719] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1720] = 32'b001111_10110_11101_0000000000000000; //['move', '$r22', '$r29']
HD[1721] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1722] = 32'b001101_00001_000000000000101101001; //['loadi', '$r1', '361']
HD[1723] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1724] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1725] = 32'b001111_10110_11110_0000000000000000; //['move', '$r22', '$r30']
HD[1726] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1727] = 32'b001101_00001_000000000000101101010; //['loadi', '$r1', '362']
HD[1728] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1729] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1730] = 32'b001111_10110_11111_0000000000000000; //['move', '$r22', '$r31']
HD[1731] = 32'b100110_00000000000000000000000000; //['flagrsrt', ' ']
HD[1732] = 32'b001101_00001_000000000000101101011; //['loadi', '$r1', '363']
HD[1733] = 32'b001110_10110_00001_0000000000000000; //['store', '$r22', '$r1']
HD[1734] = 32'b001101_11110_000000000000000010011; //['loadi', '$r30', 19]
HD[1735] = 32'b000001_00110_11000_11110_00000000000; //['add', '$r6', '$r24', '$r30']
HD[1736] = 32'b001100_00001_00110_0000000000000000; //['load', '$r1', '$r6']
HD[1737] = 32'b001101_00111_000000000000000000001; //['loadi', '$r7', '1']
HD[1738] = 32'b000001_01000_00001_00111_00000000000; //['add', '$r8', '$r1', '$r7']
HD[1739] = 32'b001101_11110_000000000000000010011; //['loadi', '$r30', 19]
HD[1740] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[1741] = 32'b001110_01000_00001_0000000000000000; //['store', '$r8', '$r1']
HD[1742] = 32'b001101_11110_000000000000000010011; //['loadi', '$r30', 19]
HD[1743] = 32'b000001_00111_11000_11110_00000000000; //['add', '$r7', '$r24', '$r30']
HD[1744] = 32'b001100_00001_00111_0000000000000000; //['load', '$r1', '$r7']
HD[1745] = 32'b001101_11110_000000000000000001101; //['loadi', '$r30', 13]
HD[1746] = 32'b000001_00111_11000_11110_00000000000; //['add', '$r7', '$r24', '$r30']
HD[1747] = 32'b001100_01000_00111_0000000000000000; //['load', '$r8', '$r7']
HD[1748] = 32'b011011_01001_00001_01000_00000000000; //['eq', '$r9', '$r1', '$r8']
HD[1749] = 32'b100010_00000_01001_0000011011011010; //['jei', '$r0', '$r9', 'L59']
HD[1750] = 32'b001101_11110_000000000000000010011; //['loadi', '$r30', 19]
HD[1751] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[1752] = 32'b001101_01001_000000000000000000000; //['loadi', '$r9', '0']
HD[1753] = 32'b001110_01001_00001_0000000000000000; //['store', '$r9', '$r1']
HD[1754] = 32'b001101_01000_000000000000000000000; //['loadi', '$r8', 0]
HD[1755] = 32'b000001_00001_11000_01000_00000000000; //['add', '$r1', '$r24', '$r8']
HD[1756] = 32'b001101_01001_000000000000000000000; //['loadi', '$r9', '0']
HD[1757] = 32'b000001_00001_00001_01001_00000000000; //['add', '$r1', '$r1', '$r9']
HD[1758] = 32'b001100_10101_00001_0000000000000000; //['load', '$r21', '$r1']
HD[1759] = 32'b001101_00001_000000000000000000000; //['loadi', '$r1', '0']
HD[1760] = 32'b011011_00011_10101_00001_00000000000; //['eq', '$r3', '$r21', '$r1']
HD[1761] = 32'b100010_00000_00011_0000011100000000; //['jei', '$r0', '$r3', 'L61']
HD[1762] = 32'b001101_00011_000000000000000000000; //['loadi', '$r3', 0]
HD[1763] = 32'b000001_00001_11000_00011_00000000000; //['add', '$r1', '$r24', '$r3']
HD[1764] = 32'b001101_00100_000000000000000000001; //['loadi', '$r4', '1']
HD[1765] = 32'b000001_00110_00001_00100_00000000000; //['add', '$r6', '$r1', '$r4']
HD[1766] = 32'b001100_00101_00110_0000000000000000; //['load', '$r5', '$r6']
HD[1767] = 32'b001101_00001_000000000000000000000; //['loadi', '$r1', '0']
HD[1768] = 32'b011011_00100_00101_00001_00000000000; //['eq', '$r4', '$r5', '$r1']
HD[1769] = 32'b100010_00000_00100_0000011100000000; //['jei', '$r0', '$r4', 'L63']
HD[1770] = 32'b001101_00100_000000000000000000000; //['loadi', '$r4', 0]
HD[1771] = 32'b000001_00001_11000_00100_00000000000; //['add', '$r1', '$r24', '$r4']
HD[1772] = 32'b001101_00101_000000000000000000010; //['loadi', '$r5', '2']
HD[1773] = 32'b000001_00111_00001_00101_00000000000; //['add', '$r7', '$r1', '$r5']
HD[1774] = 32'b001100_00110_00111_0000000000000000; //['load', '$r6', '$r7']
HD[1775] = 32'b001101_00001_000000000000000000000; //['loadi', '$r1', '0']
HD[1776] = 32'b011011_00101_00110_00001_00000000000; //['eq', '$r5', '$r6', '$r1']
HD[1777] = 32'b100010_00000_00101_0000011100000000; //['jei', '$r0', '$r5', 'L65']
HD[1778] = 32'b001101_00101_000000000000000000000; //['loadi', '$r5', 0]
HD[1779] = 32'b000001_00001_11000_00101_00000000000; //['add', '$r1', '$r24', '$r5']
HD[1780] = 32'b001101_00110_000000000000000000011; //['loadi', '$r6', '3']
HD[1781] = 32'b000001_01000_00001_00110_00000000000; //['add', '$r8', '$r1', '$r6']
HD[1782] = 32'b001100_00111_01000_0000000000000000; //['load', '$r7', '$r8']
HD[1783] = 32'b001101_00001_000000000000000000000; //['loadi', '$r1', '0']
HD[1784] = 32'b011011_00110_00111_00001_00000000000; //['eq', '$r6', '$r7', '$r1']
HD[1785] = 32'b100010_00000_00110_0000011100000000; //['jei', '$r0', '$r6', 'L67']
HD[1786] = 32'b001101_11110_000000000000000010011; //['loadi', '$r30', 19]
HD[1787] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[1788] = 32'b001101_11110_000000000000000001101; //['loadi', '$r30', 13]
HD[1789] = 32'b000001_00110_11000_11110_00000000000; //['add', '$r6', '$r24', '$r30']
HD[1790] = 32'b001100_00111_00110_0000000000000000; //['load', '$r7', '$r6']
HD[1791] = 32'b001110_00111_00001_0000000000000000; //['store', '$r7', '$r1']
HD[1792] = 32'b010000_00000_000000000000001110110; //['jmpi', 'L5']
HD[1793] = 32'b010000_00000_000000000000000000111; //['jmpi', 'L1']
HD[1794] = 32'b011001_00000000000000000000000000; // halt


//fim do programa zero





//programa um: subtraçao de duas entradas
	
		
HD[2048] = 32'b001101_00000_000000000000000000000; //['loadi', '$r0', '0']
HD[2049] = 32'b001101_11111_000000000000000000000; //['loadi', '$r31', '0']
HD[2050] = 32'b001101_11010_000000000000000000000; //['loadi', '$r26', '0']
HD[2051] = 32'b010000_00000_000000000000000000100; //['jmpi', 'main']
HD[2052] = 32'b001101_11010_000000000000000000010; //['loadi', '$r26', '2']
HD[2053] = 32'b011000_00000000000000000000000000; //['nop', ' ']
HD[2054] = 32'b101011_00000000000000000000000000; //['setprogos', ' ']
HD[2055] = 32'b011000_00000000000000000000000000; //['nop', ' ']
HD[2056] = 32'b001111_00001_11100_0000000000000000; //['move', '$r1', '$r28']
HD[2057] = 32'b001101_11110_000000000000000000000; //['loadi', '$r30', 0]
HD[2058] = 32'b000001_00010_11000_11110_00000000000; //['add', '$r2', '$r24', '$r30']
HD[2059] = 32'b001110_00001_00010_0000000000000000; //['store', '$r1', '$r2']
HD[2060] = 32'b001101_11010_000000000000000000010; //['loadi', '$r26', '2']
HD[2061] = 32'b011000_00000000000000000000000000; //['nop', ' ']
HD[2062] = 32'b101011_00000000000000000000000000; //['setprogos', ' ']
HD[2063] = 32'b011000_00000000000000000000000000; //['nop', ' ']
HD[2064] = 32'b001111_00001_11100_0000000000000000; //['move', '$r1', '$r28']
HD[2065] = 32'b001101_11110_000000000000000000001; //['loadi', '$r30', 1]
HD[2066] = 32'b000001_00010_11000_11110_00000000000; //['add', '$r2', '$r24', '$r30']
HD[2067] = 32'b001110_00001_00010_0000000000000000; //['store', '$r1', '$r2']
HD[2068] = 32'b001101_11110_000000000000000000000; //['loadi', '$r30', 0]
HD[2069] = 32'b000001_00010_11000_11110_00000000000; //['add', '$r2', '$r24', '$r30']
HD[2070] = 32'b001100_00001_00010_0000000000000000; //['load', '$r1', '$r2']
HD[2071] = 32'b001101_11110_000000000000000000001; //['loadi', '$r30', 1]
HD[2072] = 32'b000001_00010_11000_11110_00000000000; //['add', '$r2', '$r24', '$r30']
HD[2073] = 32'b001100_00011_00010_0000000000000000; //['load', '$r3', '$r2']
HD[2074] = 32'b000011_00100_00001_00011_00000000000; //['sub', '$r4', '$r1', '$r3']
HD[2075] = 32'b001101_11110_000000000000000000010; //['loadi', '$r30', 2]
HD[2076] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[2077] = 32'b001110_00100_00001_0000000000000000; //['store', '$r4', '$r1']
HD[2078] = 32'b001101_11110_000000000000000000010; //['loadi', '$r30', 2]
HD[2079] = 32'b000001_00011_11000_11110_00000000000; //['add', '$r3', '$r24', '$r30']
HD[2080] = 32'b001100_00001_00011_0000000000000000; //['load', '$r1', '$r3']
HD[2081] = 32'b001111_11001_00001_0000000000000000; //['move', '$r25', '$r1']
HD[2082] = 32'b001101_11010_000000000000000000001; //['loadi', '$r26', '1']
HD[2083] = 32'b011000_00000000000000000000000000; //['nop', ' ']
HD[2084] = 32'b101011_00000000000000000000000000; //['setprogos', ' ']
HD[2085] = 32'b011000_00000000000000000000000000; //['nop', ' ']
HD[2086] = 32'b101011_00000000000000000000000000; // setprogos

//fim programa um



//programa dois: multiplicaçao de duas entradas

HD[4096] = 32'b001101_00000_000000000000000000000; //['loadi', '$r0', '0']
HD[4097] = 32'b001101_11111_000000000000000000000; //['loadi', '$r31', '0']
HD[4098] = 32'b001101_11010_000000000000000000000; //['loadi', '$r26', '0']
HD[4099] = 32'b010000_00000_000000000000000000100; //['jmpi', 'main']
HD[4100] = 32'b001101_11010_000000000000000000010; //['loadi', '$r26', '2']
HD[4101] = 32'b011000_00000000000000000000000000; //['nop', ' ']
HD[4102] = 32'b101011_00000000000000000000000000; //['setprogos', ' ']
HD[4103] = 32'b011000_00000000000000000000000000; //['nop', ' ']
HD[4104] = 32'b001111_00001_11100_0000000000000000; //['move', '$r1', '$r28']
HD[4105] = 32'b001101_11110_000000000000000000000; //['loadi', '$r30', 0]
HD[4106] = 32'b000001_00010_11000_11110_00000000000; //['add', '$r2', '$r24', '$r30']
HD[4107] = 32'b001110_00001_00010_0000000000000000; //['store', '$r1', '$r2']
HD[4108] = 32'b001101_11010_000000000000000000010; //['loadi', '$r26', '2']
HD[4109] = 32'b011000_00000000000000000000000000; //['nop', ' ']
HD[4110] = 32'b101011_00000000000000000000000000; //['setprogos', ' ']
HD[4111] = 32'b011000_00000000000000000000000000; //['nop', ' ']
HD[4112] = 32'b001111_00001_11100_0000000000000000; //['move', '$r1', '$r28']
HD[4113] = 32'b001101_11110_000000000000000000001; //['loadi', '$r30', 1]
HD[4114] = 32'b000001_00010_11000_11110_00000000000; //['add', '$r2', '$r24', '$r30']
HD[4115] = 32'b001110_00001_00010_0000000000000000; //['store', '$r1', '$r2']
HD[4116] = 32'b001101_11110_000000000000000000000; //['loadi', '$r30', 0]
HD[4117] = 32'b000001_00010_11000_11110_00000000000; //['add', '$r2', '$r24', '$r30']
HD[4118] = 32'b001100_00001_00010_0000000000000000; //['load', '$r1', '$r2']
HD[4119] = 32'b001101_11110_000000000000000000001; //['loadi', '$r30', 1]
HD[4120] = 32'b000001_00010_11000_11110_00000000000; //['add', '$r2', '$r24', '$r30']
HD[4121] = 32'b001100_00011_00010_0000000000000000; //['load', '$r3', '$r2']
HD[4122] = 32'b000101_00100_00001_00011_00000000000; //['mult', '$r4', '$r1', '$r3']
HD[4123] = 32'b001101_11110_000000000000000000010; //['loadi', '$r30', 2]
HD[4124] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[4125] = 32'b001110_00100_00001_0000000000000000; //['store', '$r4', '$r1']
HD[4126] = 32'b001101_11110_000000000000000000010; //['loadi', '$r30', 2]
HD[4127] = 32'b000001_00011_11000_11110_00000000000; //['add', '$r3', '$r24', '$r30']
HD[4128] = 32'b001100_00001_00011_0000000000000000; //['load', '$r1', '$r3']
HD[4129] = 32'b001111_11001_00001_0000000000000000; //['move', '$r25', '$r1']
HD[4130] = 32'b001101_11010_000000000000000000001; //['loadi', '$r26', '1']
HD[4131] = 32'b011000_00000000000000000000000000; //['nop', ' ']
HD[4132] = 32'b101011_00000000000000000000000000; //['setprogos', ' ']
HD[4133] = 32'b011000_00000000000000000000000000; //['nop', ' ']
HD[4134] = 32'b101011_00000000000000000000000000; // setprogos

//fim programa dois


//programa tres: soma de dois valores

HD[6144] = 32'b001101_00000_000000000000000000000; //['loadi', '$r0', '0']
HD[6145] = 32'b001101_11111_000000000000000000000; //['loadi', '$r31', '0']
HD[6146] = 32'b001101_11010_000000000000000000000; //['loadi', '$r26', '0']
HD[6147] = 32'b010000_00000_000000000000000000100; //['jmpi', 'main']
HD[6148] = 32'b001101_11010_000000000000000000010; //['loadi', '$r26', '2']
HD[6149] = 32'b011000_00000000000000000000000000; //['nop', ' ']
HD[6150] = 32'b101011_00000000000000000000000000; //['setprogos', ' ']
HD[6151] = 32'b011000_00000000000000000000000000; //['nop', ' ']
HD[6152] = 32'b001111_00001_11100_0000000000000000; //['move', '$r1', '$r28']
HD[6153] = 32'b001101_11110_000000000000000000000; //['loadi', '$r30', 0]
HD[6154] = 32'b000001_00010_11000_11110_00000000000; //['add', '$r2', '$r24', '$r30']
HD[6155] = 32'b001110_00001_00010_0000000000000000; //['store', '$r1', '$r2']
HD[6156] = 32'b001101_11010_000000000000000000010; //['loadi', '$r26', '2']
HD[6157] = 32'b011000_00000000000000000000000000; //['nop', ' ']
HD[6158] = 32'b101011_00000000000000000000000000; //['setprogos', ' ']
HD[6159] = 32'b011000_00000000000000000000000000; //['nop', ' ']
HD[6160] = 32'b001111_00001_11100_0000000000000000; //['move', '$r1', '$r28']
HD[6161] = 32'b001101_11110_000000000000000000001; //['loadi', '$r30', 1]
HD[6162] = 32'b000001_00010_11000_11110_00000000000; //['add', '$r2', '$r24', '$r30']
HD[6163] = 32'b001110_00001_00010_0000000000000000; //['store', '$r1', '$r2']
HD[6164] = 32'b001101_11110_000000000000000000000; //['loadi', '$r30', 0]
HD[6165] = 32'b000001_00010_11000_11110_00000000000; //['add', '$r2', '$r24', '$r30']
HD[6166] = 32'b001100_00001_00010_0000000000000000; //['load', '$r1', '$r2']
HD[6167] = 32'b001101_11110_000000000000000000001; //['loadi', '$r30', 1]
HD[6168] = 32'b000001_00010_11000_11110_00000000000; //['add', '$r2', '$r24', '$r30']
HD[6169] = 32'b001100_00011_00010_0000000000000000; //['load', '$r3', '$r2']
HD[6170] = 32'b000001_00100_00001_00011_00000000000; //['add', '$r4', '$r1', '$r3']
HD[6171] = 32'b001101_11110_000000000000000000010; //['loadi', '$r30', 2]
HD[6172] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[6173] = 32'b001110_00100_00001_0000000000000000; //['store', '$r4', '$r1']
HD[6174] = 32'b001101_11110_000000000000000000010; //['loadi', '$r30', 2]
HD[6175] = 32'b000001_00011_11000_11110_00000000000; //['add', '$r3', '$r24', '$r30']
HD[6176] = 32'b001100_00001_00011_0000000000000000; //['load', '$r1', '$r3']
HD[6177] = 32'b001111_11001_00001_0000000000000000; //['move', '$r25', '$r1']
HD[6178] = 32'b001101_11010_000000000000000000001; //['loadi', '$r26', '1']
HD[6179] = 32'b011000_00000000000000000000000000; //['nop', ' ']
HD[6180] = 32'b101011_00000000000000000000000000; //['setprogos', ' ']
HD[6181] = 32'b011000_00000000000000000000000000; //['nop', ' ']
HD[6182] = 32'b101011_00000000000000000000000000; //['setprogos', ' ']

//fim programa tres



//programa quatro: fibonacci

HD[8192] = 32'b001101_00000_000000000000000000000; //['loadi', '$r0', '0']
HD[8193] = 32'b001101_11111_000000000000000000000; //['loadi', '$r31', '0']
HD[8194] = 32'b001101_11010_000000000000000000000; //['loadi', '$r26', '0']
HD[8195] = 32'b010000_00000_000000000000001010100; //['jmpi', 'main']
HD[8196] = 32'b000100_11101_11101_0000000000000001; //['subi', '$r29', '$r29', '1']
HD[8197] = 32'b100100_00001_11101_0000000000000000; //['pop', '$r1', '$r29']
HD[8198] = 32'b001101_11110_000000000000000000000; //['loadi', '$r30', 0]
HD[8199] = 32'b000001_00010_11000_11110_00000000000; //['add', '$r2', '$r24', '$r30']
HD[8200] = 32'b001110_00001_00010_0000000000000000; //['store', '$r1', '$r2']
HD[8201] = 32'b001101_11110_000000000000000000000; //['loadi', '$r30', 0]
HD[8202] = 32'b000001_00010_11000_11110_00000000000; //['add', '$r2', '$r24', '$r30']
HD[8203] = 32'b001100_00001_00010_0000000000000000; //['load', '$r1', '$r2']
HD[8204] = 32'b001101_00011_000000000000000000000; //['loadi', '$r3', '0']
HD[8205] = 32'b011110_00100_00001_00011_00000000000; //['nab', '$r4', '$r1', '$r3']
HD[8206] = 32'b100010_00000_00100_0000000000010010; //['jei', '$r0', '$r4', 'L1']
HD[8207] = 32'b001101_11100_000000000000000000000; //['loadi', '$r28', '0']
HD[8208] = 32'b010001_11111_000000000000000000000; //['jmp', '$r31']
HD[8209] = 32'b010000_00000_000000000000001010010; //['jmpi', 'L2']
HD[8210] = 32'b001101_11110_000000000000000000000; //['loadi', '$r30', 0]
HD[8211] = 32'b000001_00010_11000_11110_00000000000; //['add', '$r2', '$r24', '$r30']
HD[8212] = 32'b001100_00001_00010_0000000000000000; //['load', '$r1', '$r2']
HD[8213] = 32'b001101_00011_000000000000000000001; //['loadi', '$r3', '1']
HD[8214] = 32'b011011_00100_00001_00011_00000000000; //['eq', '$r4', '$r1', '$r3']
HD[8215] = 32'b100010_00000_00100_0000000000011011; //['jei', '$r0', '$r4', 'L3']
HD[8216] = 32'b001101_11100_000000000000000000001; //['loadi', '$r28', '1']
HD[8217] = 32'b010001_11111_000000000000000000000; //['jmp', '$r31']
HD[8218] = 32'b010000_00000_000000000000001010010; //['jmpi', 'L4']
HD[8219] = 32'b001101_11110_000000000000000000001; //['loadi', '$r30', 1]
HD[8220] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[8221] = 32'b001101_00011_000000000000000000000; //['loadi', '$r3', '0']
HD[8222] = 32'b001110_00011_00001_0000000000000000; //['store', '$r3', '$r1']
HD[8223] = 32'b001101_11110_000000000000000000010; //['loadi', '$r30', 2]
HD[8224] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[8225] = 32'b001101_00011_000000000000000000001; //['loadi', '$r3', '1']
HD[8226] = 32'b001110_00011_00001_0000000000000000; //['store', '$r3', '$r1']
HD[8227] = 32'b001101_11110_000000000000000000100; //['loadi', '$r30', 4]
HD[8228] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[8229] = 32'b001101_00011_000000000000000000001; //['loadi', '$r3', '1']
HD[8230] = 32'b001110_00011_00001_0000000000000000; //['store', '$r3', '$r1']
HD[8231] = 32'b001101_11110_000000000000000000100; //['loadi', '$r30', 4]
HD[8232] = 32'b000001_00010_11000_11110_00000000000; //['add', '$r2', '$r24', '$r30']
HD[8233] = 32'b001100_00001_00010_0000000000000000; //['load', '$r1', '$r2']
HD[8234] = 32'b001101_11110_000000000000000000000; //['loadi', '$r30', 0]
HD[8235] = 32'b000001_00010_11000_11110_00000000000; //['add', '$r2', '$r24', '$r30']
HD[8236] = 32'b001100_00011_00010_0000000000000000; //['load', '$r3', '$r2']
HD[8237] = 32'b011111_00100_00001_00011_00000000000; //['lt', '$r4', '$r1', '$r3']
HD[8238] = 32'b100010_00000_00100_0000000001001110; //['jei', '$r0', '$r4', 'L6']
HD[8239] = 32'b001101_11110_000000000000000000011; //['loadi', '$r30', 3]
HD[8240] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[8241] = 32'b001101_11110_000000000000000000010; //['loadi', '$r30', 2]
HD[8242] = 32'b000001_00011_11000_11110_00000000000; //['add', '$r3', '$r24', '$r30']
HD[8243] = 32'b001100_00100_00011_0000000000000000; //['load', '$r4', '$r3']
HD[8244] = 32'b001110_00100_00001_0000000000000000; //['store', '$r4', '$r1']
HD[8245] = 32'b001101_11110_000000000000000000010; //['loadi', '$r30', 2]
HD[8246] = 32'b000001_00011_11000_11110_00000000000; //['add', '$r3', '$r24', '$r30']
HD[8247] = 32'b001100_00001_00011_0000000000000000; //['load', '$r1', '$r3']
HD[8248] = 32'b001101_11110_000000000000000000001; //['loadi', '$r30', 1]
HD[8249] = 32'b000001_00011_11000_11110_00000000000; //['add', '$r3', '$r24', '$r30']
HD[8250] = 32'b001100_00100_00011_0000000000000000; //['load', '$r4', '$r3']
HD[8251] = 32'b000001_00101_00001_00100_00000000000; //['add', '$r5', '$r1', '$r4']
HD[8252] = 32'b001101_11110_000000000000000000010; //['loadi', '$r30', 2]
HD[8253] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[8254] = 32'b001110_00101_00001_0000000000000000; //['store', '$r5', '$r1']
HD[8255] = 32'b001101_11110_000000000000000000001; //['loadi', '$r30', 1]
HD[8256] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[8257] = 32'b001101_11110_000000000000000000011; //['loadi', '$r30', 3]
HD[8258] = 32'b000001_00100_11000_11110_00000000000; //['add', '$r4', '$r24', '$r30']
HD[8259] = 32'b001100_00101_00100_0000000000000000; //['load', '$r5', '$r4']
HD[8260] = 32'b001110_00101_00001_0000000000000000; //['store', '$r5', '$r1']
HD[8261] = 32'b001101_11110_000000000000000000100; //['loadi', '$r30', 4]
HD[8262] = 32'b000001_00100_11000_11110_00000000000; //['add', '$r4', '$r24', '$r30']
HD[8263] = 32'b001100_00001_00100_0000000000000000; //['load', '$r1', '$r4']
HD[8264] = 32'b001101_00101_000000000000000000001; //['loadi', '$r5', '1']
HD[8265] = 32'b000001_00110_00001_00101_00000000000; //['add', '$r6', '$r1', '$r5']
HD[8266] = 32'b001101_11110_000000000000000000100; //['loadi', '$r30', 4]
HD[8267] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
HD[8268] = 32'b001110_00110_00001_0000000000000000; //['store', '$r6', '$r1']
HD[8269] = 32'b010000_00000_000000000000000100111; //['jmpi', 'L5']
HD[8270] = 32'b001101_00101_000000000000000000010; //['loadi', '$r5', 2]
HD[8271] = 32'b000001_00001_11000_00101_00000000000; //['add', '$r1', '$r24', '$r5']
HD[8272] = 32'b001100_11100_00001_0000000000000000; //['load', '$r28', '$r1']
HD[8273] = 32'b010001_11111_000000000000000000000; //['jmp', '$r31']
HD[8274] = 32'b001101_11100_000000000000000000000; //['loadi', '$r28', '0']
HD[8275] = 32'b010001_11111_000000000000000000000; //['jmp', '$r31']
HD[8276] = 32'b001101_11010_000000000000000000010; //['loadi', '$r26', '2']
HD[8277] = 32'b011000_00000000000000000000000000; //['nop', ' ']
HD[8278] = 32'b101011_00000000000000000000000000; //['setprogos', ' ']
HD[8279] = 32'b011000_00000000000000000000000000; //['nop', ' ']
HD[8280] = 32'b001111_00001_11100_0000000000000000; //['move', '$r1', '$r28']
HD[8281] = 32'b001101_11110_000000000000000000101; //['loadi', '$r30', 5]
HD[8282] = 32'b000001_00010_11000_11110_00000000000; //['add', '$r2', '$r24', '$r30']
HD[8283] = 32'b001110_00001_00010_0000000000000000; //['store', '$r1', '$r2']
HD[8284] = 32'b100011_11111_11101_0000000000000000; //['push', '$r31', '$r29']
HD[8285] = 32'b000010_11101_11101_0000000000000001; //['addi', '$r29', '$r29', '1']
HD[8286] = 32'b001101_11110_000000000000000000101; //['loadi', '$r30', 5]
HD[8287] = 32'b000001_00010_11000_11110_00000000000; //['add', '$r2', '$r24', '$r30']
HD[8288] = 32'b001100_00001_00010_0000000000000000; //['load', '$r1', '$r2']
HD[8289] = 32'b100011_00001_11101_0000000000000000; //['push', '$r1', '$r29']
HD[8290] = 32'b000010_11101_11101_0000000000000001; //['addi', '$r29', '$r29', '1']
HD[8291] = 32'b100001_00000000000000000000000100; //['jal', 'fibonacci']
HD[8292] = 32'b000100_11101_11101_0000000000000001; //['subi', '$r29', '$r29', '1']
HD[8293] = 32'b100100_11111_11101_0000000000000000; //['pop', '$r31', '$r29']
HD[8294] = 32'b001111_00001_11100_0000000000000000; //['move', '$r1', '$r28']
HD[8295] = 32'b001111_11001_00001_0000000000000000; //['move', '$r25', '$r1']
HD[8296] = 32'b001101_11010_000000000000000000001; //['loadi', '$r26', '1']
HD[8297] = 32'b011000_00000000000000000000000000; //['nop', ' ']
HD[8298] = 32'b101011_00000000000000000000000000; //['setprogos', ' ']
HD[8299] = 32'b011000_00000000000000000000000000; //['nop', ' ']
HD[8300] = 32'b101011_00000000000000000000000000; //['setprogos', ' ']

//fim programa quatro



	
	end

	always @(posedge clock) begin
		
		if(write) begin // escrever dados na memória
			HD[(2048 * prog) + address] = dados_in;
		end 
		
	end
	
	
	always @(posedge clock_a) begin
		dados_out = HD[(2048 * prog) + address];
	end

endmodule