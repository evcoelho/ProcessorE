module bios(address,dados_out,clock,clock_a);
	input [31:0] address;
	input clock, clock_a;
	output reg[31:0] dados_out;
	
	reg [31:0] bios[100:0];
	
	initial begin
		//valores iniciais da bios
		
bios[0] = 32'b001101_11011_000000000000000000000; //['loadi', '$r27', '0']
bios[1] = 32'b001101_11101_000000000000000000000; //['loadi', '$r29', '0']
bios[2] = 32'b001101_11000_000000000000000000000; //['loadi', '$r24', '0']
bios[3] = 32'b001101_00000_000000000000000000000; //['loadi', '$r0', '0']
bios[4] = 32'b001101_11111_000000000000000000000; //['loadi', '$r31', '0']
bios[5] = 32'b001101_11010_000000000000000000000; //['loadi', '$r26', '0']
bios[6] = 32'b010000_00000_000000000000000000111; //['jmpi', 'main']
bios[7] = 32'b010110_11100_000000000000000000000; //['in', '$r28']
bios[8] = 32'b001111_00001_11100_0000000000000000; //['move', '$r1', '$r28']
bios[9] = 32'b001101_11110_000000000000000000001; //['loadi', '$r30', 1]
bios[10] = 32'b000001_00010_11000_11110_00000000000; //['add', '$r2', '$r24', '$r30']
bios[11] = 32'b001110_00001_00010_0000000000000000; //['store', '$r1', '$r2']
bios[12] = 32'b010110_11100_000000000000000000000; //['in', '$r28']
bios[13] = 32'b001111_00001_11100_0000000000000000; //['move', '$r1', '$r28']
bios[14] = 32'b001101_11110_000000000000000000010; //['loadi', '$r30', 2]
bios[15] = 32'b000001_00010_11000_11110_00000000000; //['add', '$r2', '$r24', '$r30']
bios[16] = 32'b001110_00001_00010_0000000000000000; //['store', '$r1', '$r2']
bios[17] = 32'b001101_11110_000000000000000000001; //['loadi', '$r30', 1]
bios[18] = 32'b000001_00010_11000_11110_00000000000; //['add', '$r2', '$r24', '$r30']
bios[19] = 32'b001100_00001_00010_0000000000000000; //['load', '$r1', '$r2']
bios[20] = 32'b001101_11110_000000000000000000010; //['loadi', '$r30', 2]
bios[21] = 32'b000001_00010_11000_11110_00000000000; //['add', '$r2', '$r24', '$r30']
bios[22] = 32'b001100_00011_00010_0000000000000000; //['load', '$r3', '$r2']
bios[23] = 32'b000001_00100_00001_00011_00000000000; //['add', '$r4', '$r1', '$r3']
bios[24] = 32'b001101_11110_000000000000000000011; //['loadi', '$r30', 3]
bios[25] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
bios[26] = 32'b001110_00100_00001_0000000000000000; //['store', '$r4', '$r1']
bios[27] = 32'b001101_11110_000000000000000000011; //['loadi', '$r30', 3]
bios[28] = 32'b000001_00011_11000_11110_00000000000; //['add', '$r3', '$r24', '$r30']
bios[29] = 32'b001100_00001_00011_0000000000000000; //['load', '$r1', '$r3']
bios[30] = 32'b010111_00001_000000000000000000000; //['out', '$r1']
bios[31] = 32'b001101_11110_000000000000000000000; //['loadi', '$r30', 0]
bios[32] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
bios[33] = 32'b001101_00100_000000000000000000000; //['loadi', '$r4', '0']
bios[34] = 32'b001110_00100_00001_0000000000000000; //['store', '$r4', '$r1']
bios[35] = 32'b001101_11110_000000000000000000000; //['loadi', '$r30', 0]
bios[36] = 32'b000001_00011_11000_11110_00000000000; //['add', '$r3', '$r24', '$r30']
bios[37] = 32'b001100_00001_00011_0000000000000000; //['load', '$r1', '$r3']
bios[38] = 32'b001101_00100_000000000011111010000; //['loadi', '$r4', '2000']
bios[39] = 32'b011111_00101_00001_00100_00000000000; //['lt', '$r5', '$r1', '$r4']
bios[40] = 32'b100010_00000_00101_0000000000111010; //['jei', '$r0', '$r5', 'L2']
bios[41] = 32'b001101_00001_000000000000000000000; //['loadi', '$r1', '0']
bios[42] = 32'b001101_11110_000000000000000000000; //['loadi', '$r30', 0]
bios[43] = 32'b000001_00100_11000_11110_00000000000; //['add', '$r4', '$r24', '$r30']
bios[44] = 32'b001100_00101_00100_0000000000000000; //['load', '$r5', '$r4']
bios[45] = 32'b001101_11110_000000000000000000000; //['loadi', '$r30', 0]
bios[46] = 32'b000001_00100_11000_11110_00000000000; //['add', '$r4', '$r24', '$r30']
bios[47] = 32'b001100_00110_00100_0000000000000000; //['load', '$r6', '$r4']
bios[48] = 32'b101010_00110_00101_00001_00000000000; //['writeosmem', '$r6', '$r5', '$r1']
bios[49] = 32'b001101_11110_000000000000000000000; //['loadi', '$r30', 0]
bios[50] = 32'b000001_00100_11000_11110_00000000000; //['add', '$r4', '$r24', '$r30']
bios[51] = 32'b001100_00001_00100_0000000000000000; //['load', '$r1', '$r4']
bios[52] = 32'b001101_00101_000000000000000000001; //['loadi', '$r5', '1']
bios[53] = 32'b000001_00110_00001_00101_00000000000; //['add', '$r6', '$r1', '$r5']
bios[54] = 32'b001101_11110_000000000000000000000; //['loadi', '$r30', 0]
bios[55] = 32'b000001_00001_11000_11110_00000000000; //['add', '$r1', '$r24', '$r30']
bios[56] = 32'b001110_00110_00001_0000000000000000; //['store', '$r6', '$r1']
bios[57] = 32'b010000_00000_000000000000000100011; //['jmpi', 'L1']
bios[58] = 32'b101110_00000000000000000000000000; // haltbios

		
		
//bios[0] = 32'b001101_00001_000000000000000000000; //['loadi', '$r1', '0'] address
//bios[1] = 32'b001101_00010_000000000000000000000; //['loadi', '$r2', '0'] prog
//bios[2] = 32'b001101_00011_000000000000000000000; //['loadi', '$r3', '0'] mem_prog
//
//bios[3] = 32'b101010_00011_00001_00010_00000000000; //['writeosmem', '$r3', '$r1', '$r2']
//bios[4] = 32'b001101_00001_000000000000000000001; //['loadi', '$r1', '1'] address
//bios[5] = 32'b001101_00011_000000000000000000001; //['loadi', '$r3', '1'] mem_prog	
//bios[6] = 32'b101010_00011_00001_00010_00000000000; //['writeosmem', '$r3', '$r1', '$r2']
//bios[7] = 32'b001101_00001_000000000000000000010; //['loadi', '$r1', '2'] address
//bios[8] = 32'b001101_00011_000000000000000000010; //['loadi', '$r3', '2'] mem_prog	
//bios[9] = 32'b101010_00011_00001_00010_00000000000; //['writeosmem', '$r3', '$r1', '$r2']
//bios[10] = 32'b101110_00000000000000000000000000; // haltBIOS
		
	end

	always @(posedge clock) begin
		
	end
	
	
	always @(posedge clock_a) begin
		dados_out = bios[address];
	end

endmodule